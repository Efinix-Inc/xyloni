`include "nt35510.vh"

module nt35510_reg
(
	input	[9:0]i_adr,
	output	[15:0]o_reg,
	output	o_dcx
);

wire	[15:0]w_reg[0:1023];
wire	[1023:0]w_dcx;

assign	w_reg[  0]	= {8'hf0, 8'h00};	assign	w_dcx[  0]	= `CMD;	assign	w_reg[  1]	= 8'h55;	assign	w_dcx[  1]	= `DAT;
assign	w_reg[  2]	= {8'hf0, 8'h01};	assign	w_dcx[  2]	= `CMD;	assign	w_reg[  3]	= 8'haa;	assign	w_dcx[  3]	= `DAT;
assign	w_reg[  4]	= {8'hf0, 8'h02};	assign	w_dcx[  4]	= `CMD;	assign	w_reg[  5]	= 8'h52;	assign	w_dcx[  5]	= `DAT;
assign	w_reg[  6]	= {8'hf0, 8'h03};	assign	w_dcx[  6]	= `CMD;	assign	w_reg[  7]	= 8'h08;	assign	w_dcx[  7]	= `DAT;
assign	w_reg[  8]	= {8'hf0, 8'h04};	assign	w_dcx[  8]	= `CMD;	assign	w_reg[  9]	= 8'h01;	assign	w_dcx[  9]	= `DAT;
assign	w_reg[ 10]	= {8'hbc, 8'h01};	assign	w_dcx[ 10]	= `CMD;	assign	w_reg[ 11]	= 8'h86;	assign	w_dcx[ 11]	= `DAT;
assign	w_reg[ 12]	= {8'hbc, 8'h02};	assign	w_dcx[ 12]	= `CMD;	assign	w_reg[ 13]	= 8'h6a;	assign	w_dcx[ 13]	= `DAT;
assign	w_reg[ 14]	= {8'hbd, 8'h01};	assign	w_dcx[ 14]	= `CMD;	assign	w_reg[ 15]	= 8'h86;	assign	w_dcx[ 15]	= `DAT;
assign	w_reg[ 16]	= {8'hbd, 8'h02};	assign	w_dcx[ 16]	= `CMD;	assign	w_reg[ 17]	= 8'h6a;	assign	w_dcx[ 17]	= `DAT;
assign	w_reg[ 18]	= {8'hbe, 8'h01};	assign	w_dcx[ 18]	= `CMD;	assign	w_reg[ 19]	= 8'h67;	assign	w_dcx[ 19]	= `DAT;
assign	w_reg[ 20]	= {8'hd1, 8'h00};	assign	w_dcx[ 20]	= `CMD;	assign	w_reg[ 21]	= 8'h00;	assign	w_dcx[ 21]	= `DAT;
assign	w_reg[ 22]	= {8'hd1, 8'h01};	assign	w_dcx[ 22]	= `CMD;	assign	w_reg[ 23]	= 8'h5d;	assign	w_dcx[ 23]	= `DAT;
assign	w_reg[ 24]	= {8'hd1, 8'h02};	assign	w_dcx[ 24]	= `CMD;	assign	w_reg[ 25]	= 8'h00;	assign	w_dcx[ 25]	= `DAT;
assign	w_reg[ 26]	= {8'hd1, 8'h03};	assign	w_dcx[ 26]	= `CMD;	assign	w_reg[ 27]	= 8'h6b;	assign	w_dcx[ 27]	= `DAT;
assign	w_reg[ 28]	= {8'hd1, 8'h04};	assign	w_dcx[ 28]	= `CMD;	assign	w_reg[ 29]	= 8'h00;	assign	w_dcx[ 29]	= `DAT;
assign	w_reg[ 30]	= {8'hd1, 8'h05};	assign	w_dcx[ 30]	= `CMD;	assign	w_reg[ 31]	= 8'h84;	assign	w_dcx[ 31]	= `DAT;
assign	w_reg[ 32]	= {8'hd1, 8'h06};	assign	w_dcx[ 32]	= `CMD;	assign	w_reg[ 33]	= 8'h00;	assign	w_dcx[ 33]	= `DAT;
assign	w_reg[ 34]	= {8'hd1, 8'h07};	assign	w_dcx[ 34]	= `CMD;	assign	w_reg[ 35]	= 8'h9c;	assign	w_dcx[ 35]	= `DAT;
assign	w_reg[ 36]	= {8'hd1, 8'h08};	assign	w_dcx[ 36]	= `CMD;	assign	w_reg[ 37]	= 8'h00;	assign	w_dcx[ 37]	= `DAT;
assign	w_reg[ 38]	= {8'hd1, 8'h09};	assign	w_dcx[ 38]	= `CMD;	assign	w_reg[ 39]	= 8'hb1;	assign	w_dcx[ 39]	= `DAT;
assign	w_reg[ 40]	= {8'hd1, 8'h0a};	assign	w_dcx[ 40]	= `CMD;	assign	w_reg[ 41]	= 8'h00;	assign	w_dcx[ 41]	= `DAT;
assign	w_reg[ 42]	= {8'hd1, 8'h0b};	assign	w_dcx[ 42]	= `CMD;	assign	w_reg[ 43]	= 8'hd9;	assign	w_dcx[ 43]	= `DAT;
assign	w_reg[ 44]	= {8'hd1, 8'h0c};	assign	w_dcx[ 44]	= `CMD;	assign	w_reg[ 45]	= 8'h00;	assign	w_dcx[ 45]	= `DAT;
assign	w_reg[ 46]	= {8'hd1, 8'h0d};	assign	w_dcx[ 46]	= `CMD;	assign	w_reg[ 47]	= 8'hfd;	assign	w_dcx[ 47]	= `DAT;
assign	w_reg[ 48]	= {8'hd1, 8'h0e};	assign	w_dcx[ 48]	= `CMD;	assign	w_reg[ 49]	= 8'h01;	assign	w_dcx[ 49]	= `DAT;
assign	w_reg[ 50]	= {8'hd1, 8'h0f};	assign	w_dcx[ 50]	= `CMD;	assign	w_reg[ 51]	= 8'h38;	assign	w_dcx[ 51]	= `DAT;
assign	w_reg[ 52]	= {8'hd1, 8'h10};	assign	w_dcx[ 52]	= `CMD;	assign	w_reg[ 53]	= 8'h01;	assign	w_dcx[ 53]	= `DAT;
assign	w_reg[ 54]	= {8'hd1, 8'h11};	assign	w_dcx[ 54]	= `CMD;	assign	w_reg[ 55]	= 8'h68;	assign	w_dcx[ 55]	= `DAT;
assign	w_reg[ 56]	= {8'hd1, 8'h12};	assign	w_dcx[ 56]	= `CMD;	assign	w_reg[ 57]	= 8'h01;	assign	w_dcx[ 57]	= `DAT;
assign	w_reg[ 58]	= {8'hd1, 8'h13};	assign	w_dcx[ 58]	= `CMD;	assign	w_reg[ 59]	= 8'hb9;	assign	w_dcx[ 59]	= `DAT;
assign	w_reg[ 60]	= {8'hd1, 8'h14};	assign	w_dcx[ 60]	= `CMD;	assign	w_reg[ 61]	= 8'h01;	assign	w_dcx[ 61]	= `DAT;
assign	w_reg[ 62]	= {8'hd1, 8'h15};	assign	w_dcx[ 62]	= `CMD;	assign	w_reg[ 63]	= 8'hfb;	assign	w_dcx[ 63]	= `DAT;
assign	w_reg[ 64]	= {8'hd1, 8'h16};	assign	w_dcx[ 64]	= `CMD;	assign	w_reg[ 65]	= 8'h02;	assign	w_dcx[ 65]	= `DAT;
assign	w_reg[ 66]	= {8'hd1, 8'h17};	assign	w_dcx[ 66]	= `CMD;	assign	w_reg[ 67]	= 8'h63;	assign	w_dcx[ 67]	= `DAT;
assign	w_reg[ 68]	= {8'hd1, 8'h18};	assign	w_dcx[ 68]	= `CMD;	assign	w_reg[ 69]	= 8'h02;	assign	w_dcx[ 69]	= `DAT;
assign	w_reg[ 70]	= {8'hd1, 8'h19};	assign	w_dcx[ 70]	= `CMD;	assign	w_reg[ 71]	= 8'hb9;	assign	w_dcx[ 71]	= `DAT;
assign	w_reg[ 72]	= {8'hd1, 8'h1a};	assign	w_dcx[ 72]	= `CMD;	assign	w_reg[ 73]	= 8'h02;	assign	w_dcx[ 73]	= `DAT;
assign	w_reg[ 74]	= {8'hd1, 8'h1b};	assign	w_dcx[ 74]	= `CMD;	assign	w_reg[ 75]	= 8'hbb;	assign	w_dcx[ 75]	= `DAT;
assign	w_reg[ 76]	= {8'hd1, 8'h1c};	assign	w_dcx[ 76]	= `CMD;	assign	w_reg[ 77]	= 8'h03;	assign	w_dcx[ 77]	= `DAT;
assign	w_reg[ 78]	= {8'hd1, 8'h1d};	assign	w_dcx[ 78]	= `CMD;	assign	w_reg[ 79]	= 8'h03;	assign	w_dcx[ 79]	= `DAT;
assign	w_reg[ 80]	= {8'hd1, 8'h1e};	assign	w_dcx[ 80]	= `CMD;	assign	w_reg[ 81]	= 8'h03;	assign	w_dcx[ 81]	= `DAT;
assign	w_reg[ 82]	= {8'hd1, 8'h1f};	assign	w_dcx[ 82]	= `CMD;	assign	w_reg[ 83]	= 8'h46;	assign	w_dcx[ 83]	= `DAT;
assign	w_reg[ 84]	= {8'hd1, 8'h20};	assign	w_dcx[ 84]	= `CMD;	assign	w_reg[ 85]	= 8'h03;	assign	w_dcx[ 85]	= `DAT;
assign	w_reg[ 86]	= {8'hd1, 8'h21};	assign	w_dcx[ 86]	= `CMD;	assign	w_reg[ 87]	= 8'h69;	assign	w_dcx[ 87]	= `DAT;
assign	w_reg[ 88]	= {8'hd1, 8'h22};	assign	w_dcx[ 88]	= `CMD;	assign	w_reg[ 89]	= 8'h03;	assign	w_dcx[ 89]	= `DAT;
assign	w_reg[ 90]	= {8'hd1, 8'h23};	assign	w_dcx[ 90]	= `CMD;	assign	w_reg[ 91]	= 8'h8f;	assign	w_dcx[ 91]	= `DAT;
assign	w_reg[ 92]	= {8'hd1, 8'h24};	assign	w_dcx[ 92]	= `CMD;	assign	w_reg[ 93]	= 8'h03;	assign	w_dcx[ 93]	= `DAT;
assign	w_reg[ 94]	= {8'hd1, 8'h25};	assign	w_dcx[ 94]	= `CMD;	assign	w_reg[ 95]	= 8'ha4;	assign	w_dcx[ 95]	= `DAT;
assign	w_reg[ 96]	= {8'hd1, 8'h26};	assign	w_dcx[ 96]	= `CMD;	assign	w_reg[ 97]	= 8'h03;	assign	w_dcx[ 97]	= `DAT;
assign	w_reg[ 98]	= {8'hd1, 8'h27};	assign	w_dcx[ 98]	= `CMD;	assign	w_reg[ 99]	= 8'hb9;	assign	w_dcx[ 99]	= `DAT;
assign	w_reg[100]	= {8'hd1, 8'h28};	assign	w_dcx[100]	= `CMD;	assign	w_reg[101]	= 8'h03;	assign	w_dcx[101]	= `DAT;
assign	w_reg[102]	= {8'hd1, 8'h29};	assign	w_dcx[102]	= `CMD;	assign	w_reg[103]	= 8'hc7;	assign	w_dcx[103]	= `DAT;
assign	w_reg[104]	= {8'hd1, 8'h2a};	assign	w_dcx[104]	= `CMD;	assign	w_reg[105]	= 8'h03;	assign	w_dcx[105]	= `DAT;
assign	w_reg[106]	= {8'hd1, 8'h2b};	assign	w_dcx[106]	= `CMD;	assign	w_reg[107]	= 8'hc9;	assign	w_dcx[107]	= `DAT;
assign	w_reg[108]	= {8'hd1, 8'h2c};	assign	w_dcx[108]	= `CMD;	assign	w_reg[109]	= 8'h03;	assign	w_dcx[109]	= `DAT;
assign	w_reg[110]	= {8'hd1, 8'h2d};	assign	w_dcx[110]	= `CMD;	assign	w_reg[111]	= 8'hcb;	assign	w_dcx[111]	= `DAT;
assign	w_reg[112]	= {8'hd1, 8'h2e};	assign	w_dcx[112]	= `CMD;	assign	w_reg[113]	= 8'h03;	assign	w_dcx[113]	= `DAT;
assign	w_reg[114]	= {8'hd1, 8'h2f};	assign	w_dcx[114]	= `CMD;	assign	w_reg[115]	= 8'hcb;	assign	w_dcx[115]	= `DAT;
assign	w_reg[116]	= {8'hd1, 8'h30};	assign	w_dcx[116]	= `CMD;	assign	w_reg[117]	= 8'h03;	assign	w_dcx[117]	= `DAT;
assign	w_reg[118]	= {8'hd1, 8'h31};	assign	w_dcx[118]	= `CMD;	assign	w_reg[119]	= 8'hcb;	assign	w_dcx[119]	= `DAT;
assign	w_reg[120]	= {8'hd1, 8'h32};	assign	w_dcx[120]	= `CMD;	assign	w_reg[121]	= 8'h03;	assign	w_dcx[121]	= `DAT;
assign	w_reg[122]	= {8'hd1, 8'h33};	assign	w_dcx[122]	= `CMD;	assign	w_reg[123]	= 8'hcc;	assign	w_dcx[123]	= `DAT;
assign	w_reg[124]	= {8'hd2, 8'h00};	assign	w_dcx[124]	= `CMD;	assign	w_reg[125]	= 8'h00;	assign	w_dcx[125]	= `DAT;
assign	w_reg[126]	= {8'hd2, 8'h01};	assign	w_dcx[126]	= `CMD;	assign	w_reg[127]	= 8'h5d;	assign	w_dcx[127]	= `DAT;
assign	w_reg[128]	= {8'hd2, 8'h02};	assign	w_dcx[128]	= `CMD;	assign	w_reg[129]	= 8'h00;	assign	w_dcx[129]	= `DAT;
assign	w_reg[130]	= {8'hd2, 8'h03};	assign	w_dcx[130]	= `CMD;	assign	w_reg[131]	= 8'h6b;	assign	w_dcx[131]	= `DAT;
assign	w_reg[132]	= {8'hd2, 8'h04};	assign	w_dcx[132]	= `CMD;	assign	w_reg[133]	= 8'h00;	assign	w_dcx[133]	= `DAT;
assign	w_reg[134]	= {8'hd2, 8'h05};	assign	w_dcx[134]	= `CMD;	assign	w_reg[135]	= 8'h84;	assign	w_dcx[135]	= `DAT;
assign	w_reg[136]	= {8'hd2, 8'h06};	assign	w_dcx[136]	= `CMD;	assign	w_reg[137]	= 8'h00;	assign	w_dcx[137]	= `DAT;
assign	w_reg[138]	= {8'hd2, 8'h07};	assign	w_dcx[138]	= `CMD;	assign	w_reg[139]	= 8'h9c;	assign	w_dcx[139]	= `DAT;
assign	w_reg[140]	= {8'hd2, 8'h08};	assign	w_dcx[140]	= `CMD;	assign	w_reg[141]	= 8'h00;	assign	w_dcx[141]	= `DAT;
assign	w_reg[142]	= {8'hd2, 8'h09};	assign	w_dcx[142]	= `CMD;	assign	w_reg[143]	= 8'hb1;	assign	w_dcx[143]	= `DAT;
assign	w_reg[144]	= {8'hd2, 8'h0a};	assign	w_dcx[144]	= `CMD;	assign	w_reg[145]	= 8'h00;	assign	w_dcx[145]	= `DAT;
assign	w_reg[146]	= {8'hd2, 8'h0b};	assign	w_dcx[146]	= `CMD;	assign	w_reg[147]	= 8'hd9;	assign	w_dcx[147]	= `DAT;
assign	w_reg[148]	= {8'hd2, 8'h0c};	assign	w_dcx[148]	= `CMD;	assign	w_reg[149]	= 8'h00;	assign	w_dcx[149]	= `DAT;
assign	w_reg[150]	= {8'hd2, 8'h0d};	assign	w_dcx[150]	= `CMD;	assign	w_reg[151]	= 8'hfd;	assign	w_dcx[151]	= `DAT;
assign	w_reg[152]	= {8'hd2, 8'h0e};	assign	w_dcx[152]	= `CMD;	assign	w_reg[153]	= 8'h01;	assign	w_dcx[153]	= `DAT;
assign	w_reg[154]	= {8'hd2, 8'h0f};	assign	w_dcx[154]	= `CMD;	assign	w_reg[155]	= 8'h38;	assign	w_dcx[155]	= `DAT;
assign	w_reg[156]	= {8'hd2, 8'h10};	assign	w_dcx[156]	= `CMD;	assign	w_reg[157]	= 8'h01;	assign	w_dcx[157]	= `DAT;
assign	w_reg[158]	= {8'hd2, 8'h11};	assign	w_dcx[158]	= `CMD;	assign	w_reg[159]	= 8'h68;	assign	w_dcx[159]	= `DAT;
assign	w_reg[160]	= {8'hd2, 8'h12};	assign	w_dcx[160]	= `CMD;	assign	w_reg[161]	= 8'h01;	assign	w_dcx[161]	= `DAT;
assign	w_reg[162]	= {8'hd2, 8'h13};	assign	w_dcx[162]	= `CMD;	assign	w_reg[163]	= 8'hb9;	assign	w_dcx[163]	= `DAT;
assign	w_reg[164]	= {8'hd2, 8'h14};	assign	w_dcx[164]	= `CMD;	assign	w_reg[165]	= 8'h01;	assign	w_dcx[165]	= `DAT;
assign	w_reg[166]	= {8'hd2, 8'h15};	assign	w_dcx[166]	= `CMD;	assign	w_reg[167]	= 8'hfb;	assign	w_dcx[167]	= `DAT;
assign	w_reg[168]	= {8'hd2, 8'h16};	assign	w_dcx[168]	= `CMD;	assign	w_reg[169]	= 8'h02;	assign	w_dcx[169]	= `DAT;
assign	w_reg[170]	= {8'hd2, 8'h17};	assign	w_dcx[170]	= `CMD;	assign	w_reg[171]	= 8'h63;	assign	w_dcx[171]	= `DAT;
assign	w_reg[172]	= {8'hd2, 8'h18};	assign	w_dcx[172]	= `CMD;	assign	w_reg[173]	= 8'h02;	assign	w_dcx[173]	= `DAT;
assign	w_reg[174]	= {8'hd2, 8'h19};	assign	w_dcx[174]	= `CMD;	assign	w_reg[175]	= 8'hb9;	assign	w_dcx[175]	= `DAT;
assign	w_reg[176]	= {8'hd2, 8'h1a};	assign	w_dcx[176]	= `CMD;	assign	w_reg[177]	= 8'h02;	assign	w_dcx[177]	= `DAT;
assign	w_reg[178]	= {8'hd2, 8'h1b};	assign	w_dcx[178]	= `CMD;	assign	w_reg[179]	= 8'hbb;	assign	w_dcx[179]	= `DAT;
assign	w_reg[180]	= {8'hd2, 8'h1c};	assign	w_dcx[180]	= `CMD;	assign	w_reg[181]	= 8'h03;	assign	w_dcx[181]	= `DAT;
assign	w_reg[182]	= {8'hd2, 8'h1d};	assign	w_dcx[182]	= `CMD;	assign	w_reg[183]	= 8'h03;	assign	w_dcx[183]	= `DAT;
assign	w_reg[184]	= {8'hd2, 8'h1e};	assign	w_dcx[184]	= `CMD;	assign	w_reg[185]	= 8'h03;	assign	w_dcx[185]	= `DAT;
assign	w_reg[186]	= {8'hd2, 8'h1f};	assign	w_dcx[186]	= `CMD;	assign	w_reg[187]	= 8'h46;	assign	w_dcx[187]	= `DAT;
assign	w_reg[188]	= {8'hd2, 8'h20};	assign	w_dcx[188]	= `CMD;	assign	w_reg[189]	= 8'h03;	assign	w_dcx[189]	= `DAT;
assign	w_reg[190]	= {8'hd2, 8'h21};	assign	w_dcx[190]	= `CMD;	assign	w_reg[191]	= 8'h69;	assign	w_dcx[191]	= `DAT;
assign	w_reg[192]	= {8'hd2, 8'h22};	assign	w_dcx[192]	= `CMD;	assign	w_reg[193]	= 8'h03;	assign	w_dcx[193]	= `DAT;
assign	w_reg[194]	= {8'hd2, 8'h23};	assign	w_dcx[194]	= `CMD;	assign	w_reg[195]	= 8'h8f;	assign	w_dcx[195]	= `DAT;
assign	w_reg[196]	= {8'hd2, 8'h24};	assign	w_dcx[196]	= `CMD;	assign	w_reg[197]	= 8'h03;	assign	w_dcx[197]	= `DAT;
assign	w_reg[198]	= {8'hd2, 8'h25};	assign	w_dcx[198]	= `CMD;	assign	w_reg[199]	= 8'ha4;	assign	w_dcx[199]	= `DAT;
assign	w_reg[200]	= {8'hd2, 8'h26};	assign	w_dcx[200]	= `CMD;	assign	w_reg[201]	= 8'h03;	assign	w_dcx[201]	= `DAT;
assign	w_reg[202]	= {8'hd2, 8'h27};	assign	w_dcx[202]	= `CMD;	assign	w_reg[203]	= 8'hb9;	assign	w_dcx[203]	= `DAT;
assign	w_reg[204]	= {8'hd2, 8'h28};	assign	w_dcx[204]	= `CMD;	assign	w_reg[205]	= 8'h03;	assign	w_dcx[205]	= `DAT;
assign	w_reg[206]	= {8'hd2, 8'h29};	assign	w_dcx[206]	= `CMD;	assign	w_reg[207]	= 8'hc7;	assign	w_dcx[207]	= `DAT;
assign	w_reg[208]	= {8'hd2, 8'h2a};	assign	w_dcx[208]	= `CMD;	assign	w_reg[209]	= 8'h03;	assign	w_dcx[209]	= `DAT;
assign	w_reg[210]	= {8'hd2, 8'h2b};	assign	w_dcx[210]	= `CMD;	assign	w_reg[211]	= 8'hc9;	assign	w_dcx[211]	= `DAT;
assign	w_reg[212]	= {8'hd2, 8'h2c};	assign	w_dcx[212]	= `CMD;	assign	w_reg[213]	= 8'h03;	assign	w_dcx[213]	= `DAT;
assign	w_reg[214]	= {8'hd2, 8'h2d};	assign	w_dcx[214]	= `CMD;	assign	w_reg[215]	= 8'hcb;	assign	w_dcx[215]	= `DAT;
assign	w_reg[216]	= {8'hd2, 8'h2e};	assign	w_dcx[216]	= `CMD;	assign	w_reg[217]	= 8'h03;	assign	w_dcx[217]	= `DAT;
assign	w_reg[218]	= {8'hd2, 8'h2f};	assign	w_dcx[218]	= `CMD;	assign	w_reg[219]	= 8'hcb;	assign	w_dcx[219]	= `DAT;
assign	w_reg[220]	= {8'hd2, 8'h30};	assign	w_dcx[220]	= `CMD;	assign	w_reg[221]	= 8'h03;	assign	w_dcx[221]	= `DAT;
assign	w_reg[222]	= {8'hd2, 8'h31};	assign	w_dcx[222]	= `CMD;	assign	w_reg[223]	= 8'hcb;	assign	w_dcx[223]	= `DAT;
assign	w_reg[224]	= {8'hd2, 8'h32};	assign	w_dcx[224]	= `CMD;	assign	w_reg[225]	= 8'h03;	assign	w_dcx[225]	= `DAT;
assign	w_reg[226]	= {8'hd2, 8'h33};	assign	w_dcx[226]	= `CMD;	assign	w_reg[227]	= 8'hcc;	assign	w_dcx[227]	= `DAT;
assign	w_reg[228]	= {8'hd3, 8'h00};	assign	w_dcx[228]	= `CMD;	assign	w_reg[229]	= 8'h00;	assign	w_dcx[229]	= `DAT;
assign	w_reg[230]	= {8'hd3, 8'h01};	assign	w_dcx[230]	= `CMD;	assign	w_reg[231]	= 8'h5d;	assign	w_dcx[231]	= `DAT;
assign	w_reg[232]	= {8'hd3, 8'h02};	assign	w_dcx[232]	= `CMD;	assign	w_reg[233]	= 8'h00;	assign	w_dcx[233]	= `DAT;
assign	w_reg[234]	= {8'hd3, 8'h03};	assign	w_dcx[234]	= `CMD;	assign	w_reg[235]	= 8'h6b;	assign	w_dcx[235]	= `DAT;
assign	w_reg[236]	= {8'hd3, 8'h04};	assign	w_dcx[236]	= `CMD;	assign	w_reg[237]	= 8'h00;	assign	w_dcx[237]	= `DAT;
assign	w_reg[238]	= {8'hd3, 8'h05};	assign	w_dcx[238]	= `CMD;	assign	w_reg[239]	= 8'h84;	assign	w_dcx[239]	= `DAT;
assign	w_reg[240]	= {8'hd3, 8'h06};	assign	w_dcx[240]	= `CMD;	assign	w_reg[241]	= 8'h00;	assign	w_dcx[241]	= `DAT;
assign	w_reg[242]	= {8'hd3, 8'h07};	assign	w_dcx[242]	= `CMD;	assign	w_reg[243]	= 8'h9c;	assign	w_dcx[243]	= `DAT;
assign	w_reg[244]	= {8'hd3, 8'h08};	assign	w_dcx[244]	= `CMD;	assign	w_reg[245]	= 8'h00;	assign	w_dcx[245]	= `DAT;
assign	w_reg[246]	= {8'hd3, 8'h09};	assign	w_dcx[246]	= `CMD;	assign	w_reg[247]	= 8'hb1;	assign	w_dcx[247]	= `DAT;
assign	w_reg[248]	= {8'hd3, 8'h0a};	assign	w_dcx[248]	= `CMD;	assign	w_reg[249]	= 8'h00;	assign	w_dcx[249]	= `DAT;
assign	w_reg[250]	= {8'hd3, 8'h0b};	assign	w_dcx[250]	= `CMD;	assign	w_reg[251]	= 8'hd9;	assign	w_dcx[251]	= `DAT;
assign	w_reg[252]	= {8'hd3, 8'h0c};	assign	w_dcx[252]	= `CMD;	assign	w_reg[253]	= 8'h00;	assign	w_dcx[253]	= `DAT;
assign	w_reg[254]	= {8'hd3, 8'h0d};	assign	w_dcx[254]	= `CMD;	assign	w_reg[255]	= 8'hfd;	assign	w_dcx[255]	= `DAT;
assign	w_reg[256]	= {8'hd3, 8'h0e};	assign	w_dcx[256]	= `CMD;	assign	w_reg[257]	= 8'h01;	assign	w_dcx[257]	= `DAT;
assign	w_reg[258]	= {8'hd3, 8'h0f};	assign	w_dcx[258]	= `CMD;	assign	w_reg[259]	= 8'h38;	assign	w_dcx[259]	= `DAT;
assign	w_reg[260]	= {8'hd3, 8'h10};	assign	w_dcx[260]	= `CMD;	assign	w_reg[261]	= 8'h01;	assign	w_dcx[261]	= `DAT;
assign	w_reg[262]	= {8'hd3, 8'h11};	assign	w_dcx[262]	= `CMD;	assign	w_reg[263]	= 8'h68;	assign	w_dcx[263]	= `DAT;
assign	w_reg[264]	= {8'hd3, 8'h12};	assign	w_dcx[264]	= `CMD;	assign	w_reg[265]	= 8'h01;	assign	w_dcx[265]	= `DAT;
assign	w_reg[266]	= {8'hd3, 8'h13};	assign	w_dcx[266]	= `CMD;	assign	w_reg[267]	= 8'hb9;	assign	w_dcx[267]	= `DAT;
assign	w_reg[268]	= {8'hd3, 8'h14};	assign	w_dcx[268]	= `CMD;	assign	w_reg[269]	= 8'h01;	assign	w_dcx[269]	= `DAT;
assign	w_reg[270]	= {8'hd3, 8'h15};	assign	w_dcx[270]	= `CMD;	assign	w_reg[271]	= 8'hfb;	assign	w_dcx[271]	= `DAT;
assign	w_reg[272]	= {8'hd3, 8'h16};	assign	w_dcx[272]	= `CMD;	assign	w_reg[273]	= 8'h02;	assign	w_dcx[273]	= `DAT;
assign	w_reg[274]	= {8'hd3, 8'h17};	assign	w_dcx[274]	= `CMD;	assign	w_reg[275]	= 8'h63;	assign	w_dcx[275]	= `DAT;
assign	w_reg[276]	= {8'hd3, 8'h18};	assign	w_dcx[276]	= `CMD;	assign	w_reg[277]	= 8'h02;	assign	w_dcx[277]	= `DAT;
assign	w_reg[278]	= {8'hd3, 8'h19};	assign	w_dcx[278]	= `CMD;	assign	w_reg[279]	= 8'hb9;	assign	w_dcx[279]	= `DAT;
assign	w_reg[280]	= {8'hd3, 8'h1a};	assign	w_dcx[280]	= `CMD;	assign	w_reg[281]	= 8'h02;	assign	w_dcx[281]	= `DAT;
assign	w_reg[282]	= {8'hd3, 8'h1b};	assign	w_dcx[282]	= `CMD;	assign	w_reg[283]	= 8'hbb;	assign	w_dcx[283]	= `DAT;
assign	w_reg[284]	= {8'hd3, 8'h1c};	assign	w_dcx[284]	= `CMD;	assign	w_reg[285]	= 8'h03;	assign	w_dcx[285]	= `DAT;
assign	w_reg[286]	= {8'hd3, 8'h1d};	assign	w_dcx[286]	= `CMD;	assign	w_reg[287]	= 8'h03;	assign	w_dcx[287]	= `DAT;
assign	w_reg[288]	= {8'hd3, 8'h1e};	assign	w_dcx[288]	= `CMD;	assign	w_reg[289]	= 8'h03;	assign	w_dcx[289]	= `DAT;
assign	w_reg[290]	= {8'hd3, 8'h1f};	assign	w_dcx[290]	= `CMD;	assign	w_reg[291]	= 8'h46;	assign	w_dcx[291]	= `DAT;
assign	w_reg[292]	= {8'hd3, 8'h20};	assign	w_dcx[292]	= `CMD;	assign	w_reg[293]	= 8'h03;	assign	w_dcx[293]	= `DAT;
assign	w_reg[294]	= {8'hd3, 8'h21};	assign	w_dcx[294]	= `CMD;	assign	w_reg[295]	= 8'h69;	assign	w_dcx[295]	= `DAT;
assign	w_reg[296]	= {8'hd3, 8'h22};	assign	w_dcx[296]	= `CMD;	assign	w_reg[297]	= 8'h03;	assign	w_dcx[297]	= `DAT;
assign	w_reg[298]	= {8'hd3, 8'h23};	assign	w_dcx[298]	= `CMD;	assign	w_reg[299]	= 8'h8f;	assign	w_dcx[299]	= `DAT;
assign	w_reg[300]	= {8'hd3, 8'h24};	assign	w_dcx[300]	= `CMD;	assign	w_reg[301]	= 8'h03;	assign	w_dcx[301]	= `DAT;
assign	w_reg[302]	= {8'hd3, 8'h25};	assign	w_dcx[302]	= `CMD;	assign	w_reg[303]	= 8'ha4;	assign	w_dcx[303]	= `DAT;
assign	w_reg[304]	= {8'hd3, 8'h26};	assign	w_dcx[304]	= `CMD;	assign	w_reg[305]	= 8'h03;	assign	w_dcx[305]	= `DAT;
assign	w_reg[306]	= {8'hd3, 8'h27};	assign	w_dcx[306]	= `CMD;	assign	w_reg[307]	= 8'hb9;	assign	w_dcx[307]	= `DAT;
assign	w_reg[308]	= {8'hd3, 8'h28};	assign	w_dcx[308]	= `CMD;	assign	w_reg[309]	= 8'h03;	assign	w_dcx[309]	= `DAT;
assign	w_reg[310]	= {8'hd3, 8'h29};	assign	w_dcx[310]	= `CMD;	assign	w_reg[311]	= 8'hc7;	assign	w_dcx[311]	= `DAT;
assign	w_reg[312]	= {8'hd3, 8'h2a};	assign	w_dcx[312]	= `CMD;	assign	w_reg[313]	= 8'h03;	assign	w_dcx[313]	= `DAT;
assign	w_reg[314]	= {8'hd3, 8'h2b};	assign	w_dcx[314]	= `CMD;	assign	w_reg[315]	= 8'hc9;	assign	w_dcx[315]	= `DAT;
assign	w_reg[316]	= {8'hd3, 8'h2c};	assign	w_dcx[316]	= `CMD;	assign	w_reg[317]	= 8'h03;	assign	w_dcx[317]	= `DAT;
assign	w_reg[318]	= {8'hd3, 8'h2d};	assign	w_dcx[318]	= `CMD;	assign	w_reg[319]	= 8'hcb;	assign	w_dcx[319]	= `DAT;
assign	w_reg[320]	= {8'hd3, 8'h2e};	assign	w_dcx[320]	= `CMD;	assign	w_reg[321]	= 8'h03;	assign	w_dcx[321]	= `DAT;
assign	w_reg[322]	= {8'hd3, 8'h2f};	assign	w_dcx[322]	= `CMD;	assign	w_reg[323]	= 8'hcb;	assign	w_dcx[323]	= `DAT;
assign	w_reg[324]	= {8'hd3, 8'h30};	assign	w_dcx[324]	= `CMD;	assign	w_reg[325]	= 8'h03;	assign	w_dcx[325]	= `DAT;
assign	w_reg[326]	= {8'hd3, 8'h31};	assign	w_dcx[326]	= `CMD;	assign	w_reg[327]	= 8'hcb;	assign	w_dcx[327]	= `DAT;
assign	w_reg[328]	= {8'hd3, 8'h32};	assign	w_dcx[328]	= `CMD;	assign	w_reg[329]	= 8'h03;	assign	w_dcx[329]	= `DAT;
assign	w_reg[330]	= {8'hd3, 8'h33};	assign	w_dcx[330]	= `CMD;	assign	w_reg[331]	= 8'hcc;	assign	w_dcx[331]	= `DAT;
assign	w_reg[332]	= {8'hd4, 8'h00};	assign	w_dcx[332]	= `CMD;	assign	w_reg[333]	= 8'h00;	assign	w_dcx[333]	= `DAT;
assign	w_reg[334]	= {8'hd4, 8'h01};	assign	w_dcx[334]	= `CMD;	assign	w_reg[335]	= 8'h5d;	assign	w_dcx[335]	= `DAT;
assign	w_reg[336]	= {8'hd4, 8'h02};	assign	w_dcx[336]	= `CMD;	assign	w_reg[337]	= 8'h00;	assign	w_dcx[337]	= `DAT;
assign	w_reg[338]	= {8'hd4, 8'h03};	assign	w_dcx[338]	= `CMD;	assign	w_reg[339]	= 8'h6b;	assign	w_dcx[339]	= `DAT;
assign	w_reg[340]	= {8'hd4, 8'h04};	assign	w_dcx[340]	= `CMD;	assign	w_reg[341]	= 8'h00;	assign	w_dcx[341]	= `DAT;
assign	w_reg[342]	= {8'hd4, 8'h05};	assign	w_dcx[342]	= `CMD;	assign	w_reg[343]	= 8'h84;	assign	w_dcx[343]	= `DAT;
assign	w_reg[344]	= {8'hd4, 8'h06};	assign	w_dcx[344]	= `CMD;	assign	w_reg[345]	= 8'h00;	assign	w_dcx[345]	= `DAT;
assign	w_reg[346]	= {8'hd4, 8'h07};	assign	w_dcx[346]	= `CMD;	assign	w_reg[347]	= 8'h9c;	assign	w_dcx[347]	= `DAT;
assign	w_reg[348]	= {8'hd4, 8'h08};	assign	w_dcx[348]	= `CMD;	assign	w_reg[349]	= 8'h00;	assign	w_dcx[349]	= `DAT;
assign	w_reg[350]	= {8'hd4, 8'h09};	assign	w_dcx[350]	= `CMD;	assign	w_reg[351]	= 8'hb1;	assign	w_dcx[351]	= `DAT;
assign	w_reg[352]	= {8'hd4, 8'h0a};	assign	w_dcx[352]	= `CMD;	assign	w_reg[353]	= 8'h00;	assign	w_dcx[353]	= `DAT;
assign	w_reg[354]	= {8'hd4, 8'h0b};	assign	w_dcx[354]	= `CMD;	assign	w_reg[355]	= 8'hd9;	assign	w_dcx[355]	= `DAT;
assign	w_reg[356]	= {8'hd4, 8'h0c};	assign	w_dcx[356]	= `CMD;	assign	w_reg[357]	= 8'h00;	assign	w_dcx[357]	= `DAT;
assign	w_reg[358]	= {8'hd4, 8'h0d};	assign	w_dcx[358]	= `CMD;	assign	w_reg[359]	= 8'hfd;	assign	w_dcx[359]	= `DAT;
assign	w_reg[360]	= {8'hd4, 8'h0e};	assign	w_dcx[360]	= `CMD;	assign	w_reg[361]	= 8'h01;	assign	w_dcx[361]	= `DAT;
assign	w_reg[362]	= {8'hd4, 8'h0f};	assign	w_dcx[362]	= `CMD;	assign	w_reg[363]	= 8'h38;	assign	w_dcx[363]	= `DAT;
assign	w_reg[364]	= {8'hd4, 8'h10};	assign	w_dcx[364]	= `CMD;	assign	w_reg[365]	= 8'h01;	assign	w_dcx[365]	= `DAT;
assign	w_reg[366]	= {8'hd4, 8'h11};	assign	w_dcx[366]	= `CMD;	assign	w_reg[367]	= 8'h68;	assign	w_dcx[367]	= `DAT;
assign	w_reg[368]	= {8'hd4, 8'h12};	assign	w_dcx[368]	= `CMD;	assign	w_reg[369]	= 8'h01;	assign	w_dcx[369]	= `DAT;
assign	w_reg[370]	= {8'hd4, 8'h13};	assign	w_dcx[370]	= `CMD;	assign	w_reg[371]	= 8'hb9;	assign	w_dcx[371]	= `DAT;
assign	w_reg[372]	= {8'hd4, 8'h14};	assign	w_dcx[372]	= `CMD;	assign	w_reg[373]	= 8'h01;	assign	w_dcx[373]	= `DAT;
assign	w_reg[374]	= {8'hd4, 8'h15};	assign	w_dcx[374]	= `CMD;	assign	w_reg[375]	= 8'hfb;	assign	w_dcx[375]	= `DAT;
assign	w_reg[376]	= {8'hd4, 8'h16};	assign	w_dcx[376]	= `CMD;	assign	w_reg[377]	= 8'h02;	assign	w_dcx[377]	= `DAT;
assign	w_reg[378]	= {8'hd4, 8'h17};	assign	w_dcx[378]	= `CMD;	assign	w_reg[379]	= 8'h63;	assign	w_dcx[379]	= `DAT;
assign	w_reg[380]	= {8'hd4, 8'h18};	assign	w_dcx[380]	= `CMD;	assign	w_reg[381]	= 8'h02;	assign	w_dcx[381]	= `DAT;
assign	w_reg[382]	= {8'hd4, 8'h19};	assign	w_dcx[382]	= `CMD;	assign	w_reg[383]	= 8'hb9;	assign	w_dcx[383]	= `DAT;
assign	w_reg[384]	= {8'hd4, 8'h1a};	assign	w_dcx[384]	= `CMD;	assign	w_reg[385]	= 8'h02;	assign	w_dcx[385]	= `DAT;
assign	w_reg[386]	= {8'hd4, 8'h1b};	assign	w_dcx[386]	= `CMD;	assign	w_reg[387]	= 8'hbb;	assign	w_dcx[387]	= `DAT;
assign	w_reg[388]	= {8'hd4, 8'h1c};	assign	w_dcx[388]	= `CMD;	assign	w_reg[389]	= 8'h03;	assign	w_dcx[389]	= `DAT;
assign	w_reg[390]	= {8'hd4, 8'h1d};	assign	w_dcx[390]	= `CMD;	assign	w_reg[391]	= 8'h03;	assign	w_dcx[391]	= `DAT;
assign	w_reg[392]	= {8'hd4, 8'h1e};	assign	w_dcx[392]	= `CMD;	assign	w_reg[393]	= 8'h03;	assign	w_dcx[393]	= `DAT;
assign	w_reg[394]	= {8'hd4, 8'h1f};	assign	w_dcx[394]	= `CMD;	assign	w_reg[395]	= 8'h46;	assign	w_dcx[395]	= `DAT;
assign	w_reg[396]	= {8'hd4, 8'h20};	assign	w_dcx[396]	= `CMD;	assign	w_reg[397]	= 8'h03;	assign	w_dcx[397]	= `DAT;
assign	w_reg[398]	= {8'hd4, 8'h21};	assign	w_dcx[398]	= `CMD;	assign	w_reg[399]	= 8'h69;	assign	w_dcx[399]	= `DAT;
assign	w_reg[400]	= {8'hd4, 8'h22};	assign	w_dcx[400]	= `CMD;	assign	w_reg[401]	= 8'h03;	assign	w_dcx[401]	= `DAT;
assign	w_reg[402]	= {8'hd4, 8'h23};	assign	w_dcx[402]	= `CMD;	assign	w_reg[403]	= 8'h8f;	assign	w_dcx[403]	= `DAT;
assign	w_reg[404]	= {8'hd4, 8'h24};	assign	w_dcx[404]	= `CMD;	assign	w_reg[405]	= 8'h03;	assign	w_dcx[405]	= `DAT;
assign	w_reg[406]	= {8'hd4, 8'h25};	assign	w_dcx[406]	= `CMD;	assign	w_reg[407]	= 8'ha4;	assign	w_dcx[407]	= `DAT;
assign	w_reg[408]	= {8'hd4, 8'h26};	assign	w_dcx[408]	= `CMD;	assign	w_reg[409]	= 8'h03;	assign	w_dcx[409]	= `DAT;
assign	w_reg[410]	= {8'hd4, 8'h27};	assign	w_dcx[410]	= `CMD;	assign	w_reg[411]	= 8'hb9;	assign	w_dcx[411]	= `DAT;
assign	w_reg[412]	= {8'hd4, 8'h28};	assign	w_dcx[412]	= `CMD;	assign	w_reg[413]	= 8'h03;	assign	w_dcx[413]	= `DAT;
assign	w_reg[414]	= {8'hd4, 8'h29};	assign	w_dcx[414]	= `CMD;	assign	w_reg[415]	= 8'hc7;	assign	w_dcx[415]	= `DAT;
assign	w_reg[416]	= {8'hd4, 8'h2a};	assign	w_dcx[416]	= `CMD;	assign	w_reg[417]	= 8'h03;	assign	w_dcx[417]	= `DAT;
assign	w_reg[418]	= {8'hd4, 8'h2b};	assign	w_dcx[418]	= `CMD;	assign	w_reg[419]	= 8'hc9;	assign	w_dcx[419]	= `DAT;
assign	w_reg[420]	= {8'hd4, 8'h2c};	assign	w_dcx[420]	= `CMD;	assign	w_reg[421]	= 8'h03;	assign	w_dcx[421]	= `DAT;
assign	w_reg[422]	= {8'hd4, 8'h2d};	assign	w_dcx[422]	= `CMD;	assign	w_reg[423]	= 8'hcb;	assign	w_dcx[423]	= `DAT;
assign	w_reg[424]	= {8'hd4, 8'h2e};	assign	w_dcx[424]	= `CMD;	assign	w_reg[425]	= 8'h03;	assign	w_dcx[425]	= `DAT;
assign	w_reg[426]	= {8'hd4, 8'h2f};	assign	w_dcx[426]	= `CMD;	assign	w_reg[427]	= 8'hcb;	assign	w_dcx[427]	= `DAT;
assign	w_reg[428]	= {8'hd4, 8'h30};	assign	w_dcx[428]	= `CMD;	assign	w_reg[429]	= 8'h03;	assign	w_dcx[429]	= `DAT;
assign	w_reg[430]	= {8'hd4, 8'h31};	assign	w_dcx[430]	= `CMD;	assign	w_reg[431]	= 8'hcb;	assign	w_dcx[431]	= `DAT;
assign	w_reg[432]	= {8'hd4, 8'h32};	assign	w_dcx[432]	= `CMD;	assign	w_reg[433]	= 8'h03;	assign	w_dcx[433]	= `DAT;
assign	w_reg[434]	= {8'hd4, 8'h33};	assign	w_dcx[434]	= `CMD;	assign	w_reg[435]	= 8'hcc;	assign	w_dcx[435]	= `DAT;
assign	w_reg[436]	= {8'hd5, 8'h00};	assign	w_dcx[436]	= `CMD;	assign	w_reg[437]	= 8'h00;	assign	w_dcx[437]	= `DAT;
assign	w_reg[438]	= {8'hd5, 8'h01};	assign	w_dcx[438]	= `CMD;	assign	w_reg[439]	= 8'h5d;	assign	w_dcx[439]	= `DAT;
assign	w_reg[440]	= {8'hd5, 8'h02};	assign	w_dcx[440]	= `CMD;	assign	w_reg[441]	= 8'h00;	assign	w_dcx[441]	= `DAT;
assign	w_reg[442]	= {8'hd5, 8'h03};	assign	w_dcx[442]	= `CMD;	assign	w_reg[443]	= 8'h6b;	assign	w_dcx[443]	= `DAT;
assign	w_reg[444]	= {8'hd5, 8'h04};	assign	w_dcx[444]	= `CMD;	assign	w_reg[445]	= 8'h00;	assign	w_dcx[445]	= `DAT;
assign	w_reg[446]	= {8'hd5, 8'h05};	assign	w_dcx[446]	= `CMD;	assign	w_reg[447]	= 8'h84;	assign	w_dcx[447]	= `DAT;
assign	w_reg[448]	= {8'hd5, 8'h06};	assign	w_dcx[448]	= `CMD;	assign	w_reg[449]	= 8'h00;	assign	w_dcx[449]	= `DAT;
assign	w_reg[450]	= {8'hd5, 8'h07};	assign	w_dcx[450]	= `CMD;	assign	w_reg[451]	= 8'h9c;	assign	w_dcx[451]	= `DAT;
assign	w_reg[452]	= {8'hd5, 8'h08};	assign	w_dcx[452]	= `CMD;	assign	w_reg[453]	= 8'h00;	assign	w_dcx[453]	= `DAT;
assign	w_reg[454]	= {8'hd5, 8'h09};	assign	w_dcx[454]	= `CMD;	assign	w_reg[455]	= 8'hb1;	assign	w_dcx[455]	= `DAT;
assign	w_reg[456]	= {8'hd5, 8'h0a};	assign	w_dcx[456]	= `CMD;	assign	w_reg[457]	= 8'h00;	assign	w_dcx[457]	= `DAT;
assign	w_reg[458]	= {8'hd5, 8'h0b};	assign	w_dcx[458]	= `CMD;	assign	w_reg[459]	= 8'hD9;	assign	w_dcx[459]	= `DAT;
assign	w_reg[460]	= {8'hd5, 8'h0c};	assign	w_dcx[460]	= `CMD;	assign	w_reg[461]	= 8'h00;	assign	w_dcx[461]	= `DAT;
assign	w_reg[462]	= {8'hd5, 8'h0d};	assign	w_dcx[462]	= `CMD;	assign	w_reg[463]	= 8'hfd;	assign	w_dcx[463]	= `DAT;
assign	w_reg[464]	= {8'hd5, 8'h0e};	assign	w_dcx[464]	= `CMD;	assign	w_reg[465]	= 8'h01;	assign	w_dcx[465]	= `DAT;
assign	w_reg[466]	= {8'hd5, 8'h0f};	assign	w_dcx[466]	= `CMD;	assign	w_reg[467]	= 8'h38;	assign	w_dcx[467]	= `DAT;
assign	w_reg[468]	= {8'hd5, 8'h10};	assign	w_dcx[468]	= `CMD;	assign	w_reg[469]	= 8'h01;	assign	w_dcx[469]	= `DAT;
assign	w_reg[470]	= {8'hd5, 8'h11};	assign	w_dcx[470]	= `CMD;	assign	w_reg[471]	= 8'h68;	assign	w_dcx[471]	= `DAT;
assign	w_reg[472]	= {8'hd5, 8'h12};	assign	w_dcx[472]	= `CMD;	assign	w_reg[473]	= 8'h01;	assign	w_dcx[473]	= `DAT;
assign	w_reg[474]	= {8'hd5, 8'h13};	assign	w_dcx[474]	= `CMD;	assign	w_reg[475]	= 8'hb9;	assign	w_dcx[475]	= `DAT;
assign	w_reg[476]	= {8'hd5, 8'h14};	assign	w_dcx[476]	= `CMD;	assign	w_reg[477]	= 8'h01;	assign	w_dcx[477]	= `DAT;
assign	w_reg[478]	= {8'hd5, 8'h15};	assign	w_dcx[478]	= `CMD;	assign	w_reg[479]	= 8'hfb;	assign	w_dcx[479]	= `DAT;
assign	w_reg[480]	= {8'hd5, 8'h16};	assign	w_dcx[480]	= `CMD;	assign	w_reg[481]	= 8'h02;	assign	w_dcx[481]	= `DAT;
assign	w_reg[482]	= {8'hd5, 8'h17};	assign	w_dcx[482]	= `CMD;	assign	w_reg[483]	= 8'h63;	assign	w_dcx[483]	= `DAT;
assign	w_reg[484]	= {8'hd5, 8'h18};	assign	w_dcx[484]	= `CMD;	assign	w_reg[485]	= 8'h02;	assign	w_dcx[485]	= `DAT;
assign	w_reg[486]	= {8'hd5, 8'h19};	assign	w_dcx[486]	= `CMD;	assign	w_reg[487]	= 8'hb9;	assign	w_dcx[487]	= `DAT;
assign	w_reg[488]	= {8'hd5, 8'h1a};	assign	w_dcx[488]	= `CMD;	assign	w_reg[489]	= 8'h02;	assign	w_dcx[489]	= `DAT;
assign	w_reg[490]	= {8'hd5, 8'h1b};	assign	w_dcx[490]	= `CMD;	assign	w_reg[491]	= 8'hbb;	assign	w_dcx[491]	= `DAT;
assign	w_reg[492]	= {8'hd5, 8'h1c};	assign	w_dcx[492]	= `CMD;	assign	w_reg[493]	= 8'h03;	assign	w_dcx[493]	= `DAT;
assign	w_reg[494]	= {8'hd5, 8'h1d};	assign	w_dcx[494]	= `CMD;	assign	w_reg[495]	= 8'h03;	assign	w_dcx[495]	= `DAT;
assign	w_reg[496]	= {8'hd5, 8'h1e};	assign	w_dcx[496]	= `CMD;	assign	w_reg[497]	= 8'h03;	assign	w_dcx[497]	= `DAT;
assign	w_reg[498]	= {8'hd5, 8'h1f};	assign	w_dcx[498]	= `CMD;	assign	w_reg[499]	= 8'h46;	assign	w_dcx[499]	= `DAT;
assign	w_reg[500]	= {8'hd5, 8'h20};	assign	w_dcx[500]	= `CMD;	assign	w_reg[501]	= 8'h03;	assign	w_dcx[501]	= `DAT;
assign	w_reg[502]	= {8'hd5, 8'h21};	assign	w_dcx[502]	= `CMD;	assign	w_reg[503]	= 8'h69;	assign	w_dcx[503]	= `DAT;
assign	w_reg[504]	= {8'hd5, 8'h22};	assign	w_dcx[504]	= `CMD;	assign	w_reg[505]	= 8'h03;	assign	w_dcx[505]	= `DAT;
assign	w_reg[506]	= {8'hd5, 8'h23};	assign	w_dcx[506]	= `CMD;	assign	w_reg[507]	= 8'h8f;	assign	w_dcx[507]	= `DAT;
assign	w_reg[508]	= {8'hd5, 8'h24};	assign	w_dcx[508]	= `CMD;	assign	w_reg[509]	= 8'h03;	assign	w_dcx[509]	= `DAT;
assign	w_reg[510]	= {8'hd5, 8'h25};	assign	w_dcx[510]	= `CMD;	assign	w_reg[511]	= 8'ha4;	assign	w_dcx[511]	= `DAT;
assign	w_reg[512]	= {8'hd5, 8'h26};	assign	w_dcx[512]	= `CMD;	assign	w_reg[513]	= 8'h03;	assign	w_dcx[513]	= `DAT;
assign	w_reg[514]	= {8'hd5, 8'h27};	assign	w_dcx[514]	= `CMD;	assign	w_reg[515]	= 8'hb9;	assign	w_dcx[515]	= `DAT;
assign	w_reg[516]	= {8'hd5, 8'h28};	assign	w_dcx[516]	= `CMD;	assign	w_reg[517]	= 8'h03;	assign	w_dcx[517]	= `DAT;
assign	w_reg[518]	= {8'hd5, 8'h29};	assign	w_dcx[518]	= `CMD;	assign	w_reg[519]	= 8'hc7;	assign	w_dcx[519]	= `DAT;
assign	w_reg[520]	= {8'hd5, 8'h2a};	assign	w_dcx[520]	= `CMD;	assign	w_reg[521]	= 8'h03;	assign	w_dcx[521]	= `DAT;
assign	w_reg[522]	= {8'hd5, 8'h2b};	assign	w_dcx[522]	= `CMD;	assign	w_reg[523]	= 8'hc9;	assign	w_dcx[523]	= `DAT;
assign	w_reg[524]	= {8'hd5, 8'h2c};	assign	w_dcx[524]	= `CMD;	assign	w_reg[525]	= 8'h03;	assign	w_dcx[525]	= `DAT;
assign	w_reg[526]	= {8'hd5, 8'h2d};	assign	w_dcx[526]	= `CMD;	assign	w_reg[527]	= 8'hcb;	assign	w_dcx[527]	= `DAT;
assign	w_reg[528]	= {8'hd5, 8'h2e};	assign	w_dcx[528]	= `CMD;	assign	w_reg[529]	= 8'h03;	assign	w_dcx[529]	= `DAT;
assign	w_reg[530]	= {8'hd5, 8'h2f};	assign	w_dcx[530]	= `CMD;	assign	w_reg[531]	= 8'hcb;	assign	w_dcx[531]	= `DAT;
assign	w_reg[532]	= {8'hd5, 8'h30};	assign	w_dcx[532]	= `CMD;	assign	w_reg[533]	= 8'h03;	assign	w_dcx[533]	= `DAT;
assign	w_reg[534]	= {8'hd5, 8'h31};	assign	w_dcx[534]	= `CMD;	assign	w_reg[535]	= 8'hcb;	assign	w_dcx[535]	= `DAT;
assign	w_reg[536]	= {8'hd5, 8'h32};	assign	w_dcx[536]	= `CMD;	assign	w_reg[537]	= 8'h03;	assign	w_dcx[537]	= `DAT;
assign	w_reg[538]	= {8'hd5, 8'h33};	assign	w_dcx[538]	= `CMD;	assign	w_reg[539]	= 8'hcc;	assign	w_dcx[539]	= `DAT;
assign	w_reg[540]	= {8'hd6, 8'h00};	assign	w_dcx[540]	= `CMD;	assign	w_reg[541]	= 8'h00;	assign	w_dcx[541]	= `DAT;
assign	w_reg[542]	= {8'hd6, 8'h01};	assign	w_dcx[542]	= `CMD;	assign	w_reg[543]	= 8'h5d;	assign	w_dcx[543]	= `DAT;
assign	w_reg[544]	= {8'hd6, 8'h02};	assign	w_dcx[544]	= `CMD;	assign	w_reg[545]	= 8'h00;	assign	w_dcx[545]	= `DAT;
assign	w_reg[546]	= {8'hd6, 8'h03};	assign	w_dcx[546]	= `CMD;	assign	w_reg[547]	= 8'h6b;	assign	w_dcx[547]	= `DAT;
assign	w_reg[548]	= {8'hd6, 8'h04};	assign	w_dcx[548]	= `CMD;	assign	w_reg[549]	= 8'h00;	assign	w_dcx[549]	= `DAT;
assign	w_reg[550]	= {8'hd6, 8'h05};	assign	w_dcx[550]	= `CMD;	assign	w_reg[551]	= 8'h84;	assign	w_dcx[551]	= `DAT;
assign	w_reg[552]	= {8'hd6, 8'h06};	assign	w_dcx[552]	= `CMD;	assign	w_reg[553]	= 8'h00;	assign	w_dcx[553]	= `DAT;
assign	w_reg[554]	= {8'hd6, 8'h07};	assign	w_dcx[554]	= `CMD;	assign	w_reg[555]	= 8'h9c;	assign	w_dcx[555]	= `DAT;
assign	w_reg[556]	= {8'hd6, 8'h08};	assign	w_dcx[556]	= `CMD;	assign	w_reg[557]	= 8'h00;	assign	w_dcx[557]	= `DAT;
assign	w_reg[558]	= {8'hd6, 8'h09};	assign	w_dcx[558]	= `CMD;	assign	w_reg[559]	= 8'hb1;	assign	w_dcx[559]	= `DAT;
assign	w_reg[560]	= {8'hd6, 8'h0a};	assign	w_dcx[560]	= `CMD;	assign	w_reg[561]	= 8'h00;	assign	w_dcx[561]	= `DAT;
assign	w_reg[562]	= {8'hd6, 8'h0b};	assign	w_dcx[562]	= `CMD;	assign	w_reg[563]	= 8'hd9;	assign	w_dcx[563]	= `DAT;
assign	w_reg[564]	= {8'hd6, 8'h0c};	assign	w_dcx[564]	= `CMD;	assign	w_reg[565]	= 8'h00;	assign	w_dcx[565]	= `DAT;
assign	w_reg[566]	= {8'hd6, 8'h0d};	assign	w_dcx[566]	= `CMD;	assign	w_reg[567]	= 8'hfd;	assign	w_dcx[567]	= `DAT;
assign	w_reg[568]	= {8'hd6, 8'h0e};	assign	w_dcx[568]	= `CMD;	assign	w_reg[569]	= 8'h01;	assign	w_dcx[569]	= `DAT;
assign	w_reg[570]	= {8'hd6, 8'h0f};	assign	w_dcx[570]	= `CMD;	assign	w_reg[571]	= 8'h38;	assign	w_dcx[571]	= `DAT;
assign	w_reg[572]	= {8'hd6, 8'h10};	assign	w_dcx[572]	= `CMD;	assign	w_reg[573]	= 8'h01;	assign	w_dcx[573]	= `DAT;
assign	w_reg[574]	= {8'hd6, 8'h11};	assign	w_dcx[574]	= `CMD;	assign	w_reg[575]	= 8'h68;	assign	w_dcx[575]	= `DAT;
assign	w_reg[576]	= {8'hd6, 8'h12};	assign	w_dcx[576]	= `CMD;	assign	w_reg[577]	= 8'h01;	assign	w_dcx[577]	= `DAT;
assign	w_reg[578]	= {8'hd6, 8'h13};	assign	w_dcx[578]	= `CMD;	assign	w_reg[579]	= 8'hb9;	assign	w_dcx[579]	= `DAT;
assign	w_reg[580]	= {8'hd6, 8'h14};	assign	w_dcx[580]	= `CMD;	assign	w_reg[581]	= 8'h01;	assign	w_dcx[581]	= `DAT;
assign	w_reg[582]	= {8'hd6, 8'h15};	assign	w_dcx[582]	= `CMD;	assign	w_reg[583]	= 8'hfb;	assign	w_dcx[583]	= `DAT;
assign	w_reg[584]	= {8'hd6, 8'h16};	assign	w_dcx[584]	= `CMD;	assign	w_reg[585]	= 8'h02;	assign	w_dcx[585]	= `DAT;
assign	w_reg[586]	= {8'hd6, 8'h17};	assign	w_dcx[586]	= `CMD;	assign	w_reg[587]	= 8'h63;	assign	w_dcx[587]	= `DAT;
assign	w_reg[588]	= {8'hd6, 8'h18};	assign	w_dcx[588]	= `CMD;	assign	w_reg[589]	= 8'h02;	assign	w_dcx[589]	= `DAT;
assign	w_reg[590]	= {8'hd6, 8'h19};	assign	w_dcx[590]	= `CMD;	assign	w_reg[591]	= 8'hb9;	assign	w_dcx[591]	= `DAT;
assign	w_reg[592]	= {8'hd6, 8'h1a};	assign	w_dcx[592]	= `CMD;	assign	w_reg[593]	= 8'h02;	assign	w_dcx[593]	= `DAT;
assign	w_reg[594]	= {8'hd6, 8'h1b};	assign	w_dcx[594]	= `CMD;	assign	w_reg[595]	= 8'hbb;	assign	w_dcx[595]	= `DAT;
assign	w_reg[596]	= {8'hd6, 8'h1c};	assign	w_dcx[596]	= `CMD;	assign	w_reg[597]	= 8'h03;	assign	w_dcx[597]	= `DAT;
assign	w_reg[598]	= {8'hd6, 8'h1d};	assign	w_dcx[598]	= `CMD;	assign	w_reg[599]	= 8'h03;	assign	w_dcx[599]	= `DAT;
assign	w_reg[600]	= {8'hd6, 8'h1e};	assign	w_dcx[600]	= `CMD;	assign	w_reg[601]	= 8'h03;	assign	w_dcx[601]	= `DAT;
assign	w_reg[602]	= {8'hd6, 8'h1f};	assign	w_dcx[602]	= `CMD;	assign	w_reg[603]	= 8'h46;	assign	w_dcx[603]	= `DAT;
assign	w_reg[604]	= {8'hd6, 8'h20};	assign	w_dcx[604]	= `CMD;	assign	w_reg[605]	= 8'h03;	assign	w_dcx[605]	= `DAT;
assign	w_reg[606]	= {8'hd6, 8'h21};	assign	w_dcx[606]	= `CMD;	assign	w_reg[607]	= 8'h69;	assign	w_dcx[607]	= `DAT;
assign	w_reg[608]	= {8'hd6, 8'h22};	assign	w_dcx[608]	= `CMD;	assign	w_reg[609]	= 8'h03;	assign	w_dcx[609]	= `DAT;
assign	w_reg[610]	= {8'hd6, 8'h23};	assign	w_dcx[610]	= `CMD;	assign	w_reg[611]	= 8'h8f;	assign	w_dcx[611]	= `DAT;
assign	w_reg[612]	= {8'hd6, 8'h24};	assign	w_dcx[612]	= `CMD;	assign	w_reg[613]	= 8'h03;	assign	w_dcx[613]	= `DAT;
assign	w_reg[614]	= {8'hd6, 8'h25};	assign	w_dcx[614]	= `CMD;	assign	w_reg[615]	= 8'ha4;	assign	w_dcx[615]	= `DAT;
assign	w_reg[616]	= {8'hd6, 8'h26};	assign	w_dcx[616]	= `CMD;	assign	w_reg[617]	= 8'h03;	assign	w_dcx[617]	= `DAT;
assign	w_reg[618]	= {8'hd6, 8'h27};	assign	w_dcx[618]	= `CMD;	assign	w_reg[619]	= 8'hb9;	assign	w_dcx[619]	= `DAT;
assign	w_reg[620]	= {8'hd6, 8'h28};	assign	w_dcx[620]	= `CMD;	assign	w_reg[621]	= 8'h03;	assign	w_dcx[621]	= `DAT;
assign	w_reg[622]	= {8'hd6, 8'h29};	assign	w_dcx[622]	= `CMD;	assign	w_reg[623]	= 8'hc7;	assign	w_dcx[623]	= `DAT;
assign	w_reg[624]	= {8'hd6, 8'h2a};	assign	w_dcx[624]	= `CMD;	assign	w_reg[625]	= 8'h03;	assign	w_dcx[625]	= `DAT;
assign	w_reg[626]	= {8'hd6, 8'h2b};	assign	w_dcx[626]	= `CMD;	assign	w_reg[627]	= 8'hc9;	assign	w_dcx[627]	= `DAT;
assign	w_reg[628]	= {8'hd6, 8'h2c};	assign	w_dcx[628]	= `CMD;	assign	w_reg[629]	= 8'h03;	assign	w_dcx[629]	= `DAT;
assign	w_reg[630]	= {8'hd6, 8'h2d};	assign	w_dcx[630]	= `CMD;	assign	w_reg[631]	= 8'hcb;	assign	w_dcx[631]	= `DAT;
assign	w_reg[632]	= {8'hd6, 8'h2e};	assign	w_dcx[632]	= `CMD;	assign	w_reg[633]	= 8'h03;	assign	w_dcx[633]	= `DAT;
assign	w_reg[634]	= {8'hd6, 8'h2f};	assign	w_dcx[634]	= `CMD;	assign	w_reg[635]	= 8'hcb;	assign	w_dcx[635]	= `DAT;
assign	w_reg[636]	= {8'hd6, 8'h30};	assign	w_dcx[636]	= `CMD;	assign	w_reg[637]	= 8'h03;	assign	w_dcx[637]	= `DAT;
assign	w_reg[638]	= {8'hd6, 8'h31};	assign	w_dcx[638]	= `CMD;	assign	w_reg[639]	= 8'hcb;	assign	w_dcx[639]	= `DAT;
assign	w_reg[640]	= {8'hd6, 8'h32};	assign	w_dcx[640]	= `CMD;	assign	w_reg[641]	= 8'h03;	assign	w_dcx[641]	= `DAT;
assign	w_reg[642]	= {8'hd6, 8'h33};	assign	w_dcx[642]	= `CMD;	assign	w_reg[643]	= 8'hcc;	assign	w_dcx[643]	= `DAT;
assign	w_reg[644]	= {8'hba, 8'h00};	assign	w_dcx[644]	= `CMD;	assign	w_reg[645]	= 8'h24;	assign	w_dcx[645]	= `DAT;
assign	w_reg[646]	= {8'hba, 8'h01};	assign	w_dcx[646]	= `CMD;	assign	w_reg[647]	= 8'h24;	assign	w_dcx[647]	= `DAT;
assign	w_reg[648]	= {8'hba, 8'h02};	assign	w_dcx[648]	= `CMD;	assign	w_reg[649]	= 8'h24;	assign	w_dcx[649]	= `DAT;
assign	w_reg[650]	= {8'hb9, 8'h00};	assign	w_dcx[650]	= `CMD;	assign	w_reg[651]	= 8'h24;	assign	w_dcx[651]	= `DAT;
assign	w_reg[652]	= {8'hb9, 8'h01};	assign	w_dcx[652]	= `CMD;	assign	w_reg[653]	= 8'h24;	assign	w_dcx[653]	= `DAT;
assign	w_reg[654]	= {8'hb9, 8'h02};	assign	w_dcx[654]	= `CMD;	assign	w_reg[655]	= 8'h24;	assign	w_dcx[655]	= `DAT;
assign	w_reg[656]	= {8'hf0, 8'h00};	assign	w_dcx[656]	= `CMD;	assign	w_reg[657]	= 8'h55;	assign	w_dcx[657]	= `DAT;
assign	w_reg[658]	= {8'hf0, 8'h01};	assign	w_dcx[658]	= `CMD;	assign	w_reg[659]	= 8'haa;	assign	w_dcx[659]	= `DAT;
assign	w_reg[660]	= {8'hf0, 8'h02};	assign	w_dcx[660]	= `CMD;	assign	w_reg[661]	= 8'h52;	assign	w_dcx[661]	= `DAT;
assign	w_reg[662]	= {8'hf0, 8'h03};	assign	w_dcx[662]	= `CMD;	assign	w_reg[663]	= 8'h08;	assign	w_dcx[663]	= `DAT;
assign	w_reg[664]	= {8'hf0, 8'h04};	assign	w_dcx[664]	= `CMD;	assign	w_reg[665]	= 8'h00;	assign	w_dcx[665]	= `DAT;
assign	w_reg[666]	= {8'hb1, 8'h00};	assign	w_dcx[666]	= `CMD;	assign	w_reg[667]	= 8'hcc;	assign	w_dcx[667]	= `DAT;
assign	w_reg[668]	= {8'hbc, 8'h00};	assign	w_dcx[668]	= `CMD;	assign	w_reg[669]	= 8'h05;	assign	w_dcx[669]	= `DAT;
assign	w_reg[670]	= {8'hbc, 8'h01};	assign	w_dcx[670]	= `CMD;	assign	w_reg[671]	= 8'h05;	assign	w_dcx[671]	= `DAT;
assign	w_reg[672]	= {8'hbc, 8'h02};	assign	w_dcx[672]	= `CMD;	assign	w_reg[673]	= 8'h05;	assign	w_dcx[673]	= `DAT;
assign	w_reg[674]	= {8'hb8, 8'h00};	assign	w_dcx[674]	= `CMD;	assign	w_reg[675]	= 8'h01;	assign	w_dcx[675]	= `DAT;
assign	w_reg[676]	= {8'hb8, 8'h01};	assign	w_dcx[676]	= `CMD;	assign	w_reg[677]	= 8'h03;	assign	w_dcx[677]	= `DAT;
assign	w_reg[678]	= {8'hb8, 8'h02};	assign	w_dcx[678]	= `CMD;	assign	w_reg[679]	= 8'h03;	assign	w_dcx[679]	= `DAT;
assign	w_reg[680]	= {8'hb8, 8'h03};	assign	w_dcx[680]	= `CMD;	assign	w_reg[681]	= 8'h03;	assign	w_dcx[681]	= `DAT;
assign	w_reg[682]	= {8'hbd, 8'h02};	assign	w_dcx[682]	= `CMD;	assign	w_reg[683]	= 8'h07;	assign	w_dcx[683]	= `DAT;
assign	w_reg[684]	= {8'hbd, 8'h03};	assign	w_dcx[684]	= `CMD;	assign	w_reg[685]	= 8'h31;	assign	w_dcx[685]	= `DAT;
assign	w_reg[686]	= {8'hbe, 8'h02};	assign	w_dcx[686]	= `CMD;	assign	w_reg[687]	= 8'h07;	assign	w_dcx[687]	= `DAT;
assign	w_reg[688]	= {8'hbe, 8'h03};	assign	w_dcx[688]	= `CMD;	assign	w_reg[689]	= 8'h31;	assign	w_dcx[689]	= `DAT;
assign	w_reg[690]	= {8'hbf, 8'h02};	assign	w_dcx[690]	= `CMD;	assign	w_reg[691]	= 8'h07;	assign	w_dcx[691]	= `DAT;
assign	w_reg[692]	= {8'hbf, 8'h03};	assign	w_dcx[692]	= `CMD;	assign	w_reg[693]	= 8'h31;	assign	w_dcx[693]	= `DAT;
assign	w_reg[694]	= {8'hff, 8'h00};	assign	w_dcx[694]	= `CMD;	assign	w_reg[695]	= 8'haa;	assign	w_dcx[695]	= `DAT;
assign	w_reg[696]	= {8'hff, 8'h01};	assign	w_dcx[696]	= `CMD;	assign	w_reg[697]	= 8'h55;	assign	w_dcx[697]	= `DAT;
assign	w_reg[698]	= {8'hff, 8'h02};	assign	w_dcx[698]	= `CMD;	assign	w_reg[699]	= 8'h25;	assign	w_dcx[699]	= `DAT;
assign	w_reg[700]	= {8'hff, 8'h03};	assign	w_dcx[700]	= `CMD;	assign	w_reg[701]	= 8'h01;	assign	w_dcx[701]	= `DAT;
assign	w_reg[702]	= {8'hf3, 8'h04};	assign	w_dcx[702]	= `CMD;	assign	w_reg[703]	= 8'h11;	assign	w_dcx[703]	= `DAT;
assign	w_reg[704]	= {8'hf3, 8'h06};	assign	w_dcx[704]	= `CMD;	assign	w_reg[705]	= 8'h10;	assign	w_dcx[705]	= `DAT;
assign	w_reg[706]	= {8'hf3, 8'h08};	assign	w_dcx[706]	= `CMD;	assign	w_reg[707]	= 8'h00;	assign	w_dcx[707]	= `DAT;

assign	w_reg[708]	= {`TEON, 8'h00};	assign	w_dcx[708]	= `CMD;	assign	w_reg[709]	= 8'h00;	assign	w_dcx[709]	= `DAT;
assign	w_reg[710]	= {`COLMOD, 8'h00};	assign	w_dcx[710]	= `CMD;	assign	w_reg[711]	= 8'h77;	assign	w_dcx[711]	= `DAT;
assign	w_reg[712]	= {`MADCTL, 8'h00};	assign	w_dcx[712]	= `CMD;	assign	w_reg[713]	= 8'h00;	assign	w_dcx[713]	= `DAT;
assign	w_reg[714]	= {`CASET, 8'h00};	assign	w_dcx[714]	= `CMD;	assign	w_reg[715]	= 8'h00;	assign	w_dcx[715]	= `DAT;	
assign	w_reg[716]	= {`CASET, 8'h01};	assign	w_dcx[716]	= `CMD;	assign	w_reg[717]	= 8'h00;	assign	w_dcx[717]	= `DAT;
assign	w_reg[718]	= {`CASET, 8'h02};	assign	w_dcx[718]	= `CMD;	assign	w_reg[719]	= 8'h01;	assign	w_dcx[719]	= `DAT;
assign	w_reg[720]	= {`CASET, 8'h03};	assign	w_dcx[720]	= `CMD;	assign	w_reg[721]	= 8'hdf;	assign	w_dcx[721]	= `DAT;
assign	w_reg[722]	= {`RASET, 8'h00};	assign	w_dcx[722]	= `CMD;	assign	w_reg[723]	= 8'h00;	assign	w_dcx[723]	= `DAT;
assign	w_reg[724]	= {`RASET, 8'h01};	assign	w_dcx[724]	= `CMD;	assign	w_reg[725]	= 8'h00;	assign	w_dcx[725]	= `DAT;
assign	w_reg[726]	= {`RASET, 8'h02};	assign	w_dcx[726]	= `CMD;	assign	w_reg[727]	= 8'h03;	assign	w_dcx[727]	= `DAT;
assign	w_reg[728]	= {`RASET, 8'h03};	assign	w_dcx[728]	= `CMD;	assign	w_reg[729]	= 8'h1f;	assign	w_dcx[729]	= `DAT;
assign	w_reg[730]	= {`SLPOUT, 8'h00};	assign	w_dcx[730]	= `CMD;	assign	w_reg[731]	= 8'h00;	assign	w_dcx[731]	= `DAT;
assign	w_reg[732]	= {`DISPON, 8'h00};	assign	w_dcx[732]	= `CMD;	assign	w_reg[733]	= 8'h00;	assign	w_dcx[733]	= `DAT;
assign	w_reg[734]	= {`RAMWR, 8'h00};	assign	w_dcx[734]	= `CMD;	assign	w_reg[735]	= 8'h00;	assign	w_dcx[735]	= `DAT;

assign	w_reg[736]	= {`DISPOFF, 8'h00};assign	w_dcx[736]	= `CMD;	assign	w_reg[737]	= 8'h00;	assign	w_dcx[737]	= `DAT;
assign	w_reg[738]	= {`SLPIN, 8'h00};	assign	w_dcx[738]	= `CMD;	assign	w_reg[739]	= 8'h00;	assign	w_dcx[739]	= `DAT;

genvar i;
generate
	for (i=740; i<1024; i=i+1)
	begin
		assign	w_reg[i] = {8'h00, 8'h00};
		assign	w_dcx[i] = 8'h00;
	end
endgenerate

assign	o_reg	= w_reg[i_adr];
assign	o_dcx	= w_dcx[i_adr];

endmodule
