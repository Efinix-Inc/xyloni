module ov5640_reg
(
	input	[9:0]i_addr,
	output	[7:0]o_data
);

wire	[(1024*8)-1:0]w_ov5640_reg;
//Initial Setting
assign	{w_ov5640_reg[(0  *24)+0*8+:8], w_ov5640_reg[(0  *24)+1*8+:8], w_ov5640_reg[(0  *24)+2*8+:8]}	= 24'h310311; // PLL Clock Select [7:2]DEBUG MODE [1]:PLL From Pad [0] DEBUG MODE
assign	{w_ov5640_reg[(1  *24)+0*8+:8], w_ov5640_reg[(1  *24)+1*8+:8], w_ov5640_reg[(1  *24)+2*8+:8]}	= 24'h300882; //SYSTEM CTROL0 System Control [7] Softwre Reset [6] Software Power Down [5:0] Debug mode
assign	{w_ov5640_reg[(2  *24)+0*8+:8], w_ov5640_reg[(2  *24)+1*8+:8], w_ov5640_reg[(2  *24)+2*8+:8]}	= 24'h300842; //SYSTEM CTROL0 System Control [7] Softwre Reset [6] Software Power Down [5:0] Debug mode
assign	{w_ov5640_reg[(3  *24)+0*8+:8], w_ov5640_reg[(3  *24)+1*8+:8], w_ov5640_reg[(3  *24)+2*8+:8]}	= 24'h310303; //SCCB SYSTEM CTRL1 PLL Clock Select [7:2]DEBUG MODE [1]:PLL From Pad [0] DEBUG MODE
assign	{w_ov5640_reg[(4  *24)+0*8+:8], w_ov5640_reg[(4  *24)+1*8+:8], w_ov5640_reg[(4  *24)+2*8+:8]}	= 24'h3017ff; //PAD OUTPUT ENABLE 01 Input/Output Control (0: input; 1: output) [7]FREX OUTPUT EN [6] VSYNC OUTPUT ENA [5] HREF OUTPUT ENA [4] PCLK OUTPUT ENA [3:0] D[9:6] OUTPUT ENA
assign	{w_ov5640_reg[(5  *24)+0*8+:8], w_ov5640_reg[(5  *24)+1*8+:8], w_ov5640_reg[(5  *24)+2*8+:8]}	= 24'h302c02; //PAD CONTROL 00 Pad Control [7:6] OUTPUT DRIVE CAPABILITY 00:1x 01:2x 10:3x 11:4x [5:2] DEBUG MODE [1]FREX ENA [0] DEBUG MODE
assign	{w_ov5640_reg[(6  *24)+0*8+:8], w_ov5640_reg[(6  *24)+1*8+:8], w_ov5640_reg[(6  *24)+2*8+:8]}	= 24'h3018ff; //PAD OUTPUT ENABLE 02 Input/Output Control (0: input; 1: output) [7:2] D[5:0] OUTPUT ENA [1] GPIO1 OUTPUT ENA [0] GPIO0 OUTPUT ENA
assign	{w_ov5640_reg[(7  *24)+0*8+:8], w_ov5640_reg[(7  *24)+1*8+:8], w_ov5640_reg[(7  *24)+2*8+:8]}	= 24'h30341A; //SC PLL CONTRL0 [7] DEBUG MODE [6:4] PLL CHARGE PUMP CONTORL [3:0] SACLE DIVIDER FOR MIPI
assign	{w_ov5640_reg[(8  *24)+0*8+:8], w_ov5640_reg[(8  *24)+1*8+:8], w_ov5640_reg[(8  *24)+2*8+:8]}	= 24'h303713; //SC PLL CONTRL3 [7:5] DEBUG MODE [4] PLL ROOT DIVIDER 0:BYPASS 1:DIV2 [3:0] PLL PRE-DIVIDER 1,2,3,4,6,8
assign	{w_ov5640_reg[(9  *24)+0*8+:8], w_ov5640_reg[(9  *24)+1*8+:8], w_ov5640_reg[(9  *24)+2*8+:8]}	= 24'h310801; //PAD OUTPUT ENABLE 02 Input/Output Control (0: input; 1: output) [7:2] D[5:0] OUTPUT ENA [1] GPIO1 OUTPUT ENA [0] GPIO0 OUTPUT ENA
assign	{w_ov5640_reg[(10 *24)+0*8+:8], w_ov5640_reg[(10 *24)+1*8+:8], w_ov5640_reg[(10 *24)+2*8+:8]}	= 24'h363036; //
assign	{w_ov5640_reg[(11 *24)+0*8+:8], w_ov5640_reg[(11 *24)+1*8+:8], w_ov5640_reg[(11 *24)+2*8+:8]}	= 24'h36310e;
assign	{w_ov5640_reg[(12 *24)+0*8+:8], w_ov5640_reg[(12 *24)+1*8+:8], w_ov5640_reg[(12 *24)+2*8+:8]}	= 24'h3632e2;
assign	{w_ov5640_reg[(13 *24)+0*8+:8], w_ov5640_reg[(13 *24)+1*8+:8], w_ov5640_reg[(13 *24)+2*8+:8]}	= 24'h363312;
assign	{w_ov5640_reg[(14 *24)+0*8+:8], w_ov5640_reg[(14 *24)+1*8+:8], w_ov5640_reg[(14 *24)+2*8+:8]}	= 24'h3621e0;
assign	{w_ov5640_reg[(15 *24)+0*8+:8], w_ov5640_reg[(15 *24)+1*8+:8], w_ov5640_reg[(15 *24)+2*8+:8]}	= 24'h3704a0;
assign	{w_ov5640_reg[(16 *24)+0*8+:8], w_ov5640_reg[(16 *24)+1*8+:8], w_ov5640_reg[(16 *24)+2*8+:8]}	= 24'h37035a;
assign	{w_ov5640_reg[(17 *24)+0*8+:8], w_ov5640_reg[(17 *24)+1*8+:8], w_ov5640_reg[(17 *24)+2*8+:8]}	= 24'h371578;
assign	{w_ov5640_reg[(18 *24)+0*8+:8], w_ov5640_reg[(18 *24)+1*8+:8], w_ov5640_reg[(18 *24)+2*8+:8]}	= 24'h371701;
assign	{w_ov5640_reg[(19 *24)+0*8+:8], w_ov5640_reg[(19 *24)+1*8+:8], w_ov5640_reg[(19 *24)+2*8+:8]}	= 24'h370b60;
assign	{w_ov5640_reg[(20 *24)+0*8+:8], w_ov5640_reg[(20 *24)+1*8+:8], w_ov5640_reg[(20 *24)+2*8+:8]}	= 24'h37051a;
assign	{w_ov5640_reg[(21 *24)+0*8+:8], w_ov5640_reg[(21 *24)+1*8+:8], w_ov5640_reg[(21 *24)+2*8+:8]}	= 24'h390502;
assign	{w_ov5640_reg[(22 *24)+0*8+:8], w_ov5640_reg[(22 *24)+1*8+:8], w_ov5640_reg[(22 *24)+2*8+:8]}	= 24'h390610;
assign	{w_ov5640_reg[(23 *24)+0*8+:8], w_ov5640_reg[(23 *24)+1*8+:8], w_ov5640_reg[(23 *24)+2*8+:8]}	= 24'h39010a;
assign	{w_ov5640_reg[(24 *24)+0*8+:8], w_ov5640_reg[(24 *24)+1*8+:8], w_ov5640_reg[(24 *24)+2*8+:8]}	= 24'h373112;
assign	{w_ov5640_reg[(25 *24)+0*8+:8], w_ov5640_reg[(25 *24)+1*8+:8], w_ov5640_reg[(25 *24)+2*8+:8]}	= 24'h360008;
assign	{w_ov5640_reg[(26 *24)+0*8+:8], w_ov5640_reg[(26 *24)+1*8+:8], w_ov5640_reg[(26 *24)+2*8+:8]}	= 24'h360133;
assign	{w_ov5640_reg[(27 *24)+0*8+:8], w_ov5640_reg[(27 *24)+1*8+:8], w_ov5640_reg[(27 *24)+2*8+:8]}	= 24'h302d60;
assign	{w_ov5640_reg[(28 *24)+0*8+:8], w_ov5640_reg[(28 *24)+1*8+:8], w_ov5640_reg[(28 *24)+2*8+:8]}	= 24'h362052;
assign	{w_ov5640_reg[(29 *24)+0*8+:8], w_ov5640_reg[(29 *24)+1*8+:8], w_ov5640_reg[(29 *24)+2*8+:8]}	= 24'h371b20;
assign	{w_ov5640_reg[(30 *24)+0*8+:8], w_ov5640_reg[(30 *24)+1*8+:8], w_ov5640_reg[(30 *24)+2*8+:8]}	= 24'h471c50;
assign	{w_ov5640_reg[(31 *24)+0*8+:8], w_ov5640_reg[(31 *24)+1*8+:8], w_ov5640_reg[(31 *24)+2*8+:8]}	= 24'h3a1343;
assign	{w_ov5640_reg[(32 *24)+0*8+:8], w_ov5640_reg[(32 *24)+1*8+:8], w_ov5640_reg[(32 *24)+2*8+:8]}	= 24'h3a1800;
assign	{w_ov5640_reg[(33 *24)+0*8+:8], w_ov5640_reg[(33 *24)+1*8+:8], w_ov5640_reg[(33 *24)+2*8+:8]}	= 24'h3a19f8;
assign	{w_ov5640_reg[(34 *24)+0*8+:8], w_ov5640_reg[(34 *24)+1*8+:8], w_ov5640_reg[(34 *24)+2*8+:8]}	= 24'h363513;
assign	{w_ov5640_reg[(35 *24)+0*8+:8], w_ov5640_reg[(35 *24)+1*8+:8], w_ov5640_reg[(35 *24)+2*8+:8]}	= 24'h363603;
assign	{w_ov5640_reg[(36 *24)+0*8+:8], w_ov5640_reg[(36 *24)+1*8+:8], w_ov5640_reg[(36 *24)+2*8+:8]}	= 24'h363440;
assign	{w_ov5640_reg[(37 *24)+0*8+:8], w_ov5640_reg[(37 *24)+1*8+:8], w_ov5640_reg[(37 *24)+2*8+:8]}	= 24'h362201;
// 50/60Hz detection
assign	{w_ov5640_reg[(38 *24)+0*8+:8], w_ov5640_reg[(38 *24)+1*8+:8], w_ov5640_reg[(38 *24)+2*8+:8]}	= 24'h3c0134;
assign	{w_ov5640_reg[(39 *24)+0*8+:8], w_ov5640_reg[(39 *24)+1*8+:8], w_ov5640_reg[(39 *24)+2*8+:8]}	= 24'h3c0428;
assign	{w_ov5640_reg[(40 *24)+0*8+:8], w_ov5640_reg[(40 *24)+1*8+:8], w_ov5640_reg[(40 *24)+2*8+:8]}	= 24'h3c0598;
assign	{w_ov5640_reg[(41 *24)+0*8+:8], w_ov5640_reg[(41 *24)+1*8+:8], w_ov5640_reg[(41 *24)+2*8+:8]}	= 24'h3c0600;
assign	{w_ov5640_reg[(42 *24)+0*8+:8], w_ov5640_reg[(42 *24)+1*8+:8], w_ov5640_reg[(42 *24)+2*8+:8]}	= 24'h3c0708;
assign	{w_ov5640_reg[(43 *24)+0*8+:8], w_ov5640_reg[(43 *24)+1*8+:8], w_ov5640_reg[(43 *24)+2*8+:8]}	= 24'h3c0800;
assign	{w_ov5640_reg[(44 *24)+0*8+:8], w_ov5640_reg[(44 *24)+1*8+:8], w_ov5640_reg[(44 *24)+2*8+:8]}	= 24'h3c091c;
assign	{w_ov5640_reg[(45 *24)+0*8+:8], w_ov5640_reg[(45 *24)+1*8+:8], w_ov5640_reg[(45 *24)+2*8+:8]}	= 24'h3c0a9c;
assign	{w_ov5640_reg[(46 *24)+0*8+:8], w_ov5640_reg[(46 *24)+1*8+:8], w_ov5640_reg[(46 *24)+2*8+:8]}	= 24'h3c0b40;
assign	{w_ov5640_reg[(47 *24)+0*8+:8], w_ov5640_reg[(47 *24)+1*8+:8], w_ov5640_reg[(47 *24)+2*8+:8]}	= 24'h381000;
assign	{w_ov5640_reg[(48 *24)+0*8+:8], w_ov5640_reg[(48 *24)+1*8+:8], w_ov5640_reg[(48 *24)+2*8+:8]}	= 24'h381110;
assign	{w_ov5640_reg[(49 *24)+0*8+:8], w_ov5640_reg[(49 *24)+1*8+:8], w_ov5640_reg[(49 *24)+2*8+:8]}	= 24'h381200;
assign	{w_ov5640_reg[(50 *24)+0*8+:8], w_ov5640_reg[(50 *24)+1*8+:8], w_ov5640_reg[(50 *24)+2*8+:8]}	= 24'h370864;
assign	{w_ov5640_reg[(51 *24)+0*8+:8], w_ov5640_reg[(51 *24)+1*8+:8], w_ov5640_reg[(51 *24)+2*8+:8]}	= 24'h400102;
assign	{w_ov5640_reg[(52 *24)+0*8+:8], w_ov5640_reg[(52 *24)+1*8+:8], w_ov5640_reg[(52 *24)+2*8+:8]}	= 24'h40051a;
assign	{w_ov5640_reg[(53 *24)+0*8+:8], w_ov5640_reg[(53 *24)+1*8+:8], w_ov5640_reg[(53 *24)+2*8+:8]}	= 24'h300000;
assign	{w_ov5640_reg[(54 *24)+0*8+:8], w_ov5640_reg[(54 *24)+1*8+:8], w_ov5640_reg[(54 *24)+2*8+:8]}	= 24'h3004ff;
assign	{w_ov5640_reg[(55 *24)+0*8+:8], w_ov5640_reg[(55 *24)+1*8+:8], w_ov5640_reg[(55 *24)+2*8+:8]}	= 24'h300e58;
assign	{w_ov5640_reg[(56 *24)+0*8+:8], w_ov5640_reg[(56 *24)+1*8+:8], w_ov5640_reg[(56 *24)+2*8+:8]}	= 24'h302e00;
assign	{w_ov5640_reg[(57 *24)+0*8+:8], w_ov5640_reg[(57 *24)+1*8+:8], w_ov5640_reg[(57 *24)+2*8+:8]}	= 24'h430060;
assign	{w_ov5640_reg[(58 *24)+0*8+:8], w_ov5640_reg[(58 *24)+1*8+:8], w_ov5640_reg[(58 *24)+2*8+:8]}	= 24'h501f01;
assign	{w_ov5640_reg[(59 *24)+0*8+:8], w_ov5640_reg[(59 *24)+1*8+:8], w_ov5640_reg[(59 *24)+2*8+:8]}	= 24'h440e00;
assign	{w_ov5640_reg[(60 *24)+0*8+:8], w_ov5640_reg[(60 *24)+1*8+:8], w_ov5640_reg[(60 *24)+2*8+:8]}	= 24'h5000a7;
// AEC target
assign	{w_ov5640_reg[(61 *24)+0*8+:8], w_ov5640_reg[(61 *24)+1*8+:8], w_ov5640_reg[(61 *24)+2*8+:8]}	= 24'h3a0f30;
assign	{w_ov5640_reg[(62 *24)+0*8+:8], w_ov5640_reg[(62 *24)+1*8+:8], w_ov5640_reg[(62 *24)+2*8+:8]}	= 24'h3a1028;
assign	{w_ov5640_reg[(63 *24)+0*8+:8], w_ov5640_reg[(63 *24)+1*8+:8], w_ov5640_reg[(63 *24)+2*8+:8]}	= 24'h3a1b30;
assign	{w_ov5640_reg[(64 *24)+0*8+:8], w_ov5640_reg[(64 *24)+1*8+:8], w_ov5640_reg[(64 *24)+2*8+:8]}	= 24'h3a1e26;
assign	{w_ov5640_reg[(65 *24)+0*8+:8], w_ov5640_reg[(65 *24)+1*8+:8], w_ov5640_reg[(65 *24)+2*8+:8]}	= 24'h3a1160;
assign	{w_ov5640_reg[(66 *24)+0*8+:8], w_ov5640_reg[(66 *24)+1*8+:8], w_ov5640_reg[(66 *24)+2*8+:8]}	= 24'h3a1f14;
// Lens correction 
assign	{w_ov5640_reg[(67 *24)+0*8+:8], w_ov5640_reg[(67 *24)+1*8+:8], w_ov5640_reg[(67 *24)+2*8+:8]}	= 24'h580023;
assign	{w_ov5640_reg[(68 *24)+0*8+:8], w_ov5640_reg[(68 *24)+1*8+:8], w_ov5640_reg[(68 *24)+2*8+:8]}	= 24'h580114;
assign	{w_ov5640_reg[(69 *24)+0*8+:8], w_ov5640_reg[(69 *24)+1*8+:8], w_ov5640_reg[(69 *24)+2*8+:8]}	= 24'h58020f;
assign	{w_ov5640_reg[(70 *24)+0*8+:8], w_ov5640_reg[(70 *24)+1*8+:8], w_ov5640_reg[(70 *24)+2*8+:8]}	= 24'h58030f;
assign	{w_ov5640_reg[(71 *24)+0*8+:8], w_ov5640_reg[(71 *24)+1*8+:8], w_ov5640_reg[(71 *24)+2*8+:8]}	= 24'h580412;
assign	{w_ov5640_reg[(72 *24)+0*8+:8], w_ov5640_reg[(72 *24)+1*8+:8], w_ov5640_reg[(72 *24)+2*8+:8]}	= 24'h580526;
assign	{w_ov5640_reg[(73 *24)+0*8+:8], w_ov5640_reg[(73 *24)+1*8+:8], w_ov5640_reg[(73 *24)+2*8+:8]}	= 24'h58060c;
assign	{w_ov5640_reg[(74 *24)+0*8+:8], w_ov5640_reg[(74 *24)+1*8+:8], w_ov5640_reg[(74 *24)+2*8+:8]}	= 24'h580708;
assign	{w_ov5640_reg[(75 *24)+0*8+:8], w_ov5640_reg[(75 *24)+1*8+:8], w_ov5640_reg[(75 *24)+2*8+:8]}	= 24'h580805;
assign	{w_ov5640_reg[(76 *24)+0*8+:8], w_ov5640_reg[(76 *24)+1*8+:8], w_ov5640_reg[(76 *24)+2*8+:8]}	= 24'h580905;
assign	{w_ov5640_reg[(77 *24)+0*8+:8], w_ov5640_reg[(77 *24)+1*8+:8], w_ov5640_reg[(77 *24)+2*8+:8]}	= 24'h580a08;
assign	{w_ov5640_reg[(78 *24)+0*8+:8], w_ov5640_reg[(78 *24)+1*8+:8], w_ov5640_reg[(78 *24)+2*8+:8]}	= 24'h580b0d;
assign	{w_ov5640_reg[(79 *24)+0*8+:8], w_ov5640_reg[(79 *24)+1*8+:8], w_ov5640_reg[(79 *24)+2*8+:8]}	= 24'h580c08;
assign	{w_ov5640_reg[(80 *24)+0*8+:8], w_ov5640_reg[(80 *24)+1*8+:8], w_ov5640_reg[(80 *24)+2*8+:8]}	= 24'h580d03;
assign	{w_ov5640_reg[(81 *24)+0*8+:8], w_ov5640_reg[(81 *24)+1*8+:8], w_ov5640_reg[(81 *24)+2*8+:8]}	= 24'h580e00;
assign	{w_ov5640_reg[(82 *24)+0*8+:8], w_ov5640_reg[(82 *24)+1*8+:8], w_ov5640_reg[(82 *24)+2*8+:8]}	= 24'h580f00;
assign	{w_ov5640_reg[(83 *24)+0*8+:8], w_ov5640_reg[(83 *24)+1*8+:8], w_ov5640_reg[(83 *24)+2*8+:8]}	= 24'h581003;
assign	{w_ov5640_reg[(84 *24)+0*8+:8], w_ov5640_reg[(84 *24)+1*8+:8], w_ov5640_reg[(84 *24)+2*8+:8]}	= 24'h581109;
assign	{w_ov5640_reg[(85 *24)+0*8+:8], w_ov5640_reg[(85 *24)+1*8+:8], w_ov5640_reg[(85 *24)+2*8+:8]}	= 24'h581207;
assign	{w_ov5640_reg[(86 *24)+0*8+:8], w_ov5640_reg[(86 *24)+1*8+:8], w_ov5640_reg[(86 *24)+2*8+:8]}	= 24'h581303;
assign	{w_ov5640_reg[(87 *24)+0*8+:8], w_ov5640_reg[(87 *24)+1*8+:8], w_ov5640_reg[(87 *24)+2*8+:8]}	= 24'h581400;
assign	{w_ov5640_reg[(88 *24)+0*8+:8], w_ov5640_reg[(88 *24)+1*8+:8], w_ov5640_reg[(88 *24)+2*8+:8]}	= 24'h581501;
assign	{w_ov5640_reg[(89 *24)+0*8+:8], w_ov5640_reg[(89 *24)+1*8+:8], w_ov5640_reg[(89 *24)+2*8+:8]}	= 24'h581603;
assign	{w_ov5640_reg[(90 *24)+0*8+:8], w_ov5640_reg[(90 *24)+1*8+:8], w_ov5640_reg[(90 *24)+2*8+:8]}	= 24'h581708;
assign	{w_ov5640_reg[(91 *24)+0*8+:8], w_ov5640_reg[(91 *24)+1*8+:8], w_ov5640_reg[(91 *24)+2*8+:8]}	= 24'h58180d;
assign	{w_ov5640_reg[(92 *24)+0*8+:8], w_ov5640_reg[(92 *24)+1*8+:8], w_ov5640_reg[(92 *24)+2*8+:8]}	= 24'h581908;
assign	{w_ov5640_reg[(93 *24)+0*8+:8], w_ov5640_reg[(93 *24)+1*8+:8], w_ov5640_reg[(93 *24)+2*8+:8]}	= 24'h581a05;
assign	{w_ov5640_reg[(94 *24)+0*8+:8], w_ov5640_reg[(94 *24)+1*8+:8], w_ov5640_reg[(94 *24)+2*8+:8]}	= 24'h581b06;
assign	{w_ov5640_reg[(95 *24)+0*8+:8], w_ov5640_reg[(95 *24)+1*8+:8], w_ov5640_reg[(95 *24)+2*8+:8]}	= 24'h581c08;
assign	{w_ov5640_reg[(96 *24)+0*8+:8], w_ov5640_reg[(96 *24)+1*8+:8], w_ov5640_reg[(96 *24)+2*8+:8]}	= 24'h581d0e;
assign	{w_ov5640_reg[(97 *24)+0*8+:8], w_ov5640_reg[(97 *24)+1*8+:8], w_ov5640_reg[(97 *24)+2*8+:8]}	= 24'h581e29;
assign	{w_ov5640_reg[(98 *24)+0*8+:8], w_ov5640_reg[(98 *24)+1*8+:8], w_ov5640_reg[(98 *24)+2*8+:8]}	= 24'h581f17;
assign	{w_ov5640_reg[(99 *24)+0*8+:8], w_ov5640_reg[(99 *24)+1*8+:8], w_ov5640_reg[(99 *24)+2*8+:8]}	= 24'h582011;
assign	{w_ov5640_reg[(100*24)+0*8+:8], w_ov5640_reg[(100*24)+1*8+:8], w_ov5640_reg[(100*24)+2*8+:8]}	= 24'h582111;
assign	{w_ov5640_reg[(101*24)+0*8+:8], w_ov5640_reg[(101*24)+1*8+:8], w_ov5640_reg[(101*24)+2*8+:8]}	= 24'h582215;
assign	{w_ov5640_reg[(102*24)+0*8+:8], w_ov5640_reg[(102*24)+1*8+:8], w_ov5640_reg[(102*24)+2*8+:8]}	= 24'h582328;
assign	{w_ov5640_reg[(103*24)+0*8+:8], w_ov5640_reg[(103*24)+1*8+:8], w_ov5640_reg[(103*24)+2*8+:8]}	= 24'h582446;
assign	{w_ov5640_reg[(104*24)+0*8+:8], w_ov5640_reg[(104*24)+1*8+:8], w_ov5640_reg[(104*24)+2*8+:8]}	= 24'h582526;
assign	{w_ov5640_reg[(105*24)+0*8+:8], w_ov5640_reg[(105*24)+1*8+:8], w_ov5640_reg[(105*24)+2*8+:8]}	= 24'h582608;
assign	{w_ov5640_reg[(106*24)+0*8+:8], w_ov5640_reg[(106*24)+1*8+:8], w_ov5640_reg[(106*24)+2*8+:8]}	= 24'h582726;
assign	{w_ov5640_reg[(107*24)+0*8+:8], w_ov5640_reg[(107*24)+1*8+:8], w_ov5640_reg[(107*24)+2*8+:8]}	= 24'h582864;
assign	{w_ov5640_reg[(108*24)+0*8+:8], w_ov5640_reg[(108*24)+1*8+:8], w_ov5640_reg[(108*24)+2*8+:8]}	= 24'h582926;
assign	{w_ov5640_reg[(109*24)+0*8+:8], w_ov5640_reg[(109*24)+1*8+:8], w_ov5640_reg[(109*24)+2*8+:8]}	= 24'h582a24;
assign	{w_ov5640_reg[(110*24)+0*8+:8], w_ov5640_reg[(110*24)+1*8+:8], w_ov5640_reg[(110*24)+2*8+:8]}	= 24'h582b22;
assign	{w_ov5640_reg[(111*24)+0*8+:8], w_ov5640_reg[(111*24)+1*8+:8], w_ov5640_reg[(111*24)+2*8+:8]}	= 24'h582c24;
assign	{w_ov5640_reg[(112*24)+0*8+:8], w_ov5640_reg[(112*24)+1*8+:8], w_ov5640_reg[(112*24)+2*8+:8]}	= 24'h582d24;
assign	{w_ov5640_reg[(113*24)+0*8+:8], w_ov5640_reg[(113*24)+1*8+:8], w_ov5640_reg[(113*24)+2*8+:8]}	= 24'h582e06;
assign	{w_ov5640_reg[(114*24)+0*8+:8], w_ov5640_reg[(114*24)+1*8+:8], w_ov5640_reg[(114*24)+2*8+:8]}	= 24'h582f22;
assign	{w_ov5640_reg[(115*24)+0*8+:8], w_ov5640_reg[(115*24)+1*8+:8], w_ov5640_reg[(115*24)+2*8+:8]}	= 24'h583040;
assign	{w_ov5640_reg[(116*24)+0*8+:8], w_ov5640_reg[(116*24)+1*8+:8], w_ov5640_reg[(116*24)+2*8+:8]}	= 24'h583142;
assign	{w_ov5640_reg[(117*24)+0*8+:8], w_ov5640_reg[(117*24)+1*8+:8], w_ov5640_reg[(117*24)+2*8+:8]}	= 24'h583224;
assign	{w_ov5640_reg[(118*24)+0*8+:8], w_ov5640_reg[(118*24)+1*8+:8], w_ov5640_reg[(118*24)+2*8+:8]}	= 24'h583326;
assign	{w_ov5640_reg[(119*24)+0*8+:8], w_ov5640_reg[(119*24)+1*8+:8], w_ov5640_reg[(119*24)+2*8+:8]}	= 24'h583424;
assign	{w_ov5640_reg[(120*24)+0*8+:8], w_ov5640_reg[(120*24)+1*8+:8], w_ov5640_reg[(120*24)+2*8+:8]}	= 24'h583522;
assign	{w_ov5640_reg[(121*24)+0*8+:8], w_ov5640_reg[(121*24)+1*8+:8], w_ov5640_reg[(121*24)+2*8+:8]}	= 24'h583622;
assign	{w_ov5640_reg[(122*24)+0*8+:8], w_ov5640_reg[(122*24)+1*8+:8], w_ov5640_reg[(122*24)+2*8+:8]}	= 24'h583726;
assign	{w_ov5640_reg[(123*24)+0*8+:8], w_ov5640_reg[(123*24)+1*8+:8], w_ov5640_reg[(123*24)+2*8+:8]}	= 24'h583844;
assign	{w_ov5640_reg[(124*24)+0*8+:8], w_ov5640_reg[(124*24)+1*8+:8], w_ov5640_reg[(124*24)+2*8+:8]}	= 24'h583924;
assign	{w_ov5640_reg[(125*24)+0*8+:8], w_ov5640_reg[(125*24)+1*8+:8], w_ov5640_reg[(125*24)+2*8+:8]}	= 24'h583a26;
assign	{w_ov5640_reg[(126*24)+0*8+:8], w_ov5640_reg[(126*24)+1*8+:8], w_ov5640_reg[(126*24)+2*8+:8]}	= 24'h583b28;
assign	{w_ov5640_reg[(127*24)+0*8+:8], w_ov5640_reg[(127*24)+1*8+:8], w_ov5640_reg[(127*24)+2*8+:8]}	= 24'h583c42;
assign	{w_ov5640_reg[(128*24)+0*8+:8], w_ov5640_reg[(128*24)+1*8+:8], w_ov5640_reg[(128*24)+2*8+:8]}	= 24'h583dce;
//AWB
assign	{w_ov5640_reg[(129*24)+0*8+:8], w_ov5640_reg[(129*24)+1*8+:8], w_ov5640_reg[(129*24)+2*8+:8]}	= 24'h5180ff;
assign	{w_ov5640_reg[(130*24)+0*8+:8], w_ov5640_reg[(130*24)+1*8+:8], w_ov5640_reg[(130*24)+2*8+:8]}	= 24'h5181f2;
assign	{w_ov5640_reg[(131*24)+0*8+:8], w_ov5640_reg[(131*24)+1*8+:8], w_ov5640_reg[(131*24)+2*8+:8]}	= 24'h518200;
assign	{w_ov5640_reg[(132*24)+0*8+:8], w_ov5640_reg[(132*24)+1*8+:8], w_ov5640_reg[(132*24)+2*8+:8]}	= 24'h518314;
assign	{w_ov5640_reg[(133*24)+0*8+:8], w_ov5640_reg[(133*24)+1*8+:8], w_ov5640_reg[(133*24)+2*8+:8]}	= 24'h518425;
assign	{w_ov5640_reg[(134*24)+0*8+:8], w_ov5640_reg[(134*24)+1*8+:8], w_ov5640_reg[(134*24)+2*8+:8]}	= 24'h518524;
assign	{w_ov5640_reg[(135*24)+0*8+:8], w_ov5640_reg[(135*24)+1*8+:8], w_ov5640_reg[(135*24)+2*8+:8]}	= 24'h518609;
assign	{w_ov5640_reg[(136*24)+0*8+:8], w_ov5640_reg[(136*24)+1*8+:8], w_ov5640_reg[(136*24)+2*8+:8]}	= 24'h518709;
assign	{w_ov5640_reg[(137*24)+0*8+:8], w_ov5640_reg[(137*24)+1*8+:8], w_ov5640_reg[(137*24)+2*8+:8]}	= 24'h518809;
assign	{w_ov5640_reg[(138*24)+0*8+:8], w_ov5640_reg[(138*24)+1*8+:8], w_ov5640_reg[(138*24)+2*8+:8]}	= 24'h518975;
assign	{w_ov5640_reg[(139*24)+0*8+:8], w_ov5640_reg[(139*24)+1*8+:8], w_ov5640_reg[(139*24)+2*8+:8]}	= 24'h518a54;
assign	{w_ov5640_reg[(140*24)+0*8+:8], w_ov5640_reg[(140*24)+1*8+:8], w_ov5640_reg[(140*24)+2*8+:8]}	= 24'h518be0;
assign	{w_ov5640_reg[(141*24)+0*8+:8], w_ov5640_reg[(141*24)+1*8+:8], w_ov5640_reg[(141*24)+2*8+:8]}	= 24'h518cb2;
assign	{w_ov5640_reg[(142*24)+0*8+:8], w_ov5640_reg[(142*24)+1*8+:8], w_ov5640_reg[(142*24)+2*8+:8]}	= 24'h518d42;
assign	{w_ov5640_reg[(143*24)+0*8+:8], w_ov5640_reg[(143*24)+1*8+:8], w_ov5640_reg[(143*24)+2*8+:8]}	= 24'h518e3d;
assign	{w_ov5640_reg[(144*24)+0*8+:8], w_ov5640_reg[(144*24)+1*8+:8], w_ov5640_reg[(144*24)+2*8+:8]}	= 24'h518f56;
assign	{w_ov5640_reg[(145*24)+0*8+:8], w_ov5640_reg[(145*24)+1*8+:8], w_ov5640_reg[(145*24)+2*8+:8]}	= 24'h519046;
assign	{w_ov5640_reg[(146*24)+0*8+:8], w_ov5640_reg[(146*24)+1*8+:8], w_ov5640_reg[(146*24)+2*8+:8]}	= 24'h5191f8;
assign	{w_ov5640_reg[(147*24)+0*8+:8], w_ov5640_reg[(147*24)+1*8+:8], w_ov5640_reg[(147*24)+2*8+:8]}	= 24'h519204;
assign	{w_ov5640_reg[(148*24)+0*8+:8], w_ov5640_reg[(148*24)+1*8+:8], w_ov5640_reg[(148*24)+2*8+:8]}	= 24'h5193f0;
assign	{w_ov5640_reg[(149*24)+0*8+:8], w_ov5640_reg[(149*24)+1*8+:8], w_ov5640_reg[(149*24)+2*8+:8]}	= 24'h519470;
assign	{w_ov5640_reg[(150*24)+0*8+:8], w_ov5640_reg[(150*24)+1*8+:8], w_ov5640_reg[(150*24)+2*8+:8]}	= 24'h5195f0;
assign	{w_ov5640_reg[(151*24)+0*8+:8], w_ov5640_reg[(151*24)+1*8+:8], w_ov5640_reg[(151*24)+2*8+:8]}	= 24'h519603;
assign	{w_ov5640_reg[(152*24)+0*8+:8], w_ov5640_reg[(152*24)+1*8+:8], w_ov5640_reg[(152*24)+2*8+:8]}	= 24'h519701;
assign	{w_ov5640_reg[(153*24)+0*8+:8], w_ov5640_reg[(153*24)+1*8+:8], w_ov5640_reg[(153*24)+2*8+:8]}	= 24'h519804;
assign	{w_ov5640_reg[(154*24)+0*8+:8], w_ov5640_reg[(154*24)+1*8+:8], w_ov5640_reg[(154*24)+2*8+:8]}	= 24'h519912;
assign	{w_ov5640_reg[(155*24)+0*8+:8], w_ov5640_reg[(155*24)+1*8+:8], w_ov5640_reg[(155*24)+2*8+:8]}	= 24'h519a04;
assign	{w_ov5640_reg[(156*24)+0*8+:8], w_ov5640_reg[(156*24)+1*8+:8], w_ov5640_reg[(156*24)+2*8+:8]}	= 24'h519b00;
assign	{w_ov5640_reg[(157*24)+0*8+:8], w_ov5640_reg[(157*24)+1*8+:8], w_ov5640_reg[(157*24)+2*8+:8]}	= 24'h519c06;
assign	{w_ov5640_reg[(158*24)+0*8+:8], w_ov5640_reg[(158*24)+1*8+:8], w_ov5640_reg[(158*24)+2*8+:8]}	= 24'h519d82;
assign	{w_ov5640_reg[(159*24)+0*8+:8], w_ov5640_reg[(159*24)+1*8+:8], w_ov5640_reg[(159*24)+2*8+:8]}	= 24'h519e38;
// Gamma
assign	{w_ov5640_reg[(160*24)+0*8+:8], w_ov5640_reg[(160*24)+1*8+:8], w_ov5640_reg[(160*24)+2*8+:8]}	= 24'h548001;
assign	{w_ov5640_reg[(161*24)+0*8+:8], w_ov5640_reg[(161*24)+1*8+:8], w_ov5640_reg[(161*24)+2*8+:8]}	= 24'h548108;
assign	{w_ov5640_reg[(162*24)+0*8+:8], w_ov5640_reg[(162*24)+1*8+:8], w_ov5640_reg[(162*24)+2*8+:8]}	= 24'h548214;
assign	{w_ov5640_reg[(163*24)+0*8+:8], w_ov5640_reg[(163*24)+1*8+:8], w_ov5640_reg[(163*24)+2*8+:8]}	= 24'h548328;
assign	{w_ov5640_reg[(164*24)+0*8+:8], w_ov5640_reg[(164*24)+1*8+:8], w_ov5640_reg[(164*24)+2*8+:8]}	= 24'h548451;
assign	{w_ov5640_reg[(165*24)+0*8+:8], w_ov5640_reg[(165*24)+1*8+:8], w_ov5640_reg[(165*24)+2*8+:8]}	= 24'h548565;
assign	{w_ov5640_reg[(166*24)+0*8+:8], w_ov5640_reg[(166*24)+1*8+:8], w_ov5640_reg[(166*24)+2*8+:8]}	= 24'h548671;
assign	{w_ov5640_reg[(167*24)+0*8+:8], w_ov5640_reg[(167*24)+1*8+:8], w_ov5640_reg[(167*24)+2*8+:8]}	= 24'h54877d;
assign	{w_ov5640_reg[(168*24)+0*8+:8], w_ov5640_reg[(168*24)+1*8+:8], w_ov5640_reg[(168*24)+2*8+:8]}	= 24'h548887;
assign	{w_ov5640_reg[(169*24)+0*8+:8], w_ov5640_reg[(169*24)+1*8+:8], w_ov5640_reg[(169*24)+2*8+:8]}	= 24'h548991;
assign	{w_ov5640_reg[(170*24)+0*8+:8], w_ov5640_reg[(170*24)+1*8+:8], w_ov5640_reg[(170*24)+2*8+:8]}	= 24'h548a9a;
assign	{w_ov5640_reg[(171*24)+0*8+:8], w_ov5640_reg[(171*24)+1*8+:8], w_ov5640_reg[(171*24)+2*8+:8]}	= 24'h548baa;
assign	{w_ov5640_reg[(172*24)+0*8+:8], w_ov5640_reg[(172*24)+1*8+:8], w_ov5640_reg[(172*24)+2*8+:8]}	= 24'h548cb8;
assign	{w_ov5640_reg[(173*24)+0*8+:8], w_ov5640_reg[(173*24)+1*8+:8], w_ov5640_reg[(173*24)+2*8+:8]}	= 24'h548dcd;
assign	{w_ov5640_reg[(174*24)+0*8+:8], w_ov5640_reg[(174*24)+1*8+:8], w_ov5640_reg[(174*24)+2*8+:8]}	= 24'h548edd;
assign	{w_ov5640_reg[(175*24)+0*8+:8], w_ov5640_reg[(175*24)+1*8+:8], w_ov5640_reg[(175*24)+2*8+:8]}	= 24'h548fea;
assign	{w_ov5640_reg[(176*24)+0*8+:8], w_ov5640_reg[(176*24)+1*8+:8], w_ov5640_reg[(176*24)+2*8+:8]}	= 24'h54901d;
// color matrix
assign	{w_ov5640_reg[(177*24)+0*8+:8], w_ov5640_reg[(177*24)+1*8+:8], w_ov5640_reg[(177*24)+2*8+:8]}	= 24'h53811e;
assign	{w_ov5640_reg[(178*24)+0*8+:8], w_ov5640_reg[(178*24)+1*8+:8], w_ov5640_reg[(178*24)+2*8+:8]}	= 24'h53825b;
assign	{w_ov5640_reg[(179*24)+0*8+:8], w_ov5640_reg[(179*24)+1*8+:8], w_ov5640_reg[(179*24)+2*8+:8]}	= 24'h538308;
assign	{w_ov5640_reg[(180*24)+0*8+:8], w_ov5640_reg[(180*24)+1*8+:8], w_ov5640_reg[(180*24)+2*8+:8]}	= 24'h53840a;
assign	{w_ov5640_reg[(181*24)+0*8+:8], w_ov5640_reg[(181*24)+1*8+:8], w_ov5640_reg[(181*24)+2*8+:8]}	= 24'h53857e;
assign	{w_ov5640_reg[(182*24)+0*8+:8], w_ov5640_reg[(182*24)+1*8+:8], w_ov5640_reg[(182*24)+2*8+:8]}	= 24'h538688;
assign	{w_ov5640_reg[(183*24)+0*8+:8], w_ov5640_reg[(183*24)+1*8+:8], w_ov5640_reg[(183*24)+2*8+:8]}	= 24'h53877c;
assign	{w_ov5640_reg[(184*24)+0*8+:8], w_ov5640_reg[(184*24)+1*8+:8], w_ov5640_reg[(184*24)+2*8+:8]}	= 24'h53886c;
assign	{w_ov5640_reg[(185*24)+0*8+:8], w_ov5640_reg[(185*24)+1*8+:8], w_ov5640_reg[(185*24)+2*8+:8]}	= 24'h538910;
assign	{w_ov5640_reg[(186*24)+0*8+:8], w_ov5640_reg[(186*24)+1*8+:8], w_ov5640_reg[(186*24)+2*8+:8]}	= 24'h538a01;
assign	{w_ov5640_reg[(187*24)+0*8+:8], w_ov5640_reg[(187*24)+1*8+:8], w_ov5640_reg[(187*24)+2*8+:8]}	= 24'h538b98;
// UV adjsut
assign	{w_ov5640_reg[(188*24)+0*8+:8], w_ov5640_reg[(188*24)+1*8+:8], w_ov5640_reg[(188*24)+2*8+:8]}	= 24'h558006;
assign	{w_ov5640_reg[(189*24)+0*8+:8], w_ov5640_reg[(189*24)+1*8+:8], w_ov5640_reg[(189*24)+2*8+:8]}	= 24'h558340;
assign	{w_ov5640_reg[(190*24)+0*8+:8], w_ov5640_reg[(190*24)+1*8+:8], w_ov5640_reg[(190*24)+2*8+:8]}	= 24'h558410;
assign	{w_ov5640_reg[(191*24)+0*8+:8], w_ov5640_reg[(191*24)+1*8+:8], w_ov5640_reg[(191*24)+2*8+:8]}	= 24'h558910;
assign	{w_ov5640_reg[(192*24)+0*8+:8], w_ov5640_reg[(192*24)+1*8+:8], w_ov5640_reg[(192*24)+2*8+:8]}	= 24'h558a00;
assign	{w_ov5640_reg[(193*24)+0*8+:8], w_ov5640_reg[(193*24)+1*8+:8], w_ov5640_reg[(193*24)+2*8+:8]}	= 24'h558bf8;
assign	{w_ov5640_reg[(194*24)+0*8+:8], w_ov5640_reg[(194*24)+1*8+:8], w_ov5640_reg[(194*24)+2*8+:8]}	= 24'h501d40;
// CIP
assign	{w_ov5640_reg[(195*24)+0*8+:8], w_ov5640_reg[(195*24)+1*8+:8], w_ov5640_reg[(195*24)+2*8+:8]}	= 24'h530008;
assign	{w_ov5640_reg[(196*24)+0*8+:8], w_ov5640_reg[(196*24)+1*8+:8], w_ov5640_reg[(196*24)+2*8+:8]}	= 24'h530130;
assign	{w_ov5640_reg[(197*24)+0*8+:8], w_ov5640_reg[(197*24)+1*8+:8], w_ov5640_reg[(197*24)+2*8+:8]}	= 24'h530210;
assign	{w_ov5640_reg[(198*24)+0*8+:8], w_ov5640_reg[(198*24)+1*8+:8], w_ov5640_reg[(198*24)+2*8+:8]}	= 24'h530300;
assign	{w_ov5640_reg[(199*24)+0*8+:8], w_ov5640_reg[(199*24)+1*8+:8], w_ov5640_reg[(199*24)+2*8+:8]}	= 24'h530408;
assign	{w_ov5640_reg[(200*24)+0*8+:8], w_ov5640_reg[(200*24)+1*8+:8], w_ov5640_reg[(200*24)+2*8+:8]}	= 24'h530530;
assign	{w_ov5640_reg[(201*24)+0*8+:8], w_ov5640_reg[(201*24)+1*8+:8], w_ov5640_reg[(201*24)+2*8+:8]}	= 24'h530608;
assign	{w_ov5640_reg[(202*24)+0*8+:8], w_ov5640_reg[(202*24)+1*8+:8], w_ov5640_reg[(202*24)+2*8+:8]}	= 24'h530716;
assign	{w_ov5640_reg[(203*24)+0*8+:8], w_ov5640_reg[(203*24)+1*8+:8], w_ov5640_reg[(203*24)+2*8+:8]}	= 24'h530908;
assign	{w_ov5640_reg[(204*24)+0*8+:8], w_ov5640_reg[(204*24)+1*8+:8], w_ov5640_reg[(204*24)+2*8+:8]}	= 24'h530a30;
assign	{w_ov5640_reg[(205*24)+0*8+:8], w_ov5640_reg[(205*24)+1*8+:8], w_ov5640_reg[(205*24)+2*8+:8]}	= 24'h530b04;
assign	{w_ov5640_reg[(206*24)+0*8+:8], w_ov5640_reg[(206*24)+1*8+:8], w_ov5640_reg[(206*24)+2*8+:8]}	= 24'h530c06;
assign	{w_ov5640_reg[(207*24)+0*8+:8], w_ov5640_reg[(207*24)+1*8+:8], w_ov5640_reg[(207*24)+2*8+:8]}	= 24'h502500;
assign	{w_ov5640_reg[(208*24)+0*8+:8], w_ov5640_reg[(208*24)+1*8+:8], w_ov5640_reg[(208*24)+2*8+:8]}	= 24'h300802;

//720p
assign	{w_ov5640_reg[(209*24)+0*8+:8], w_ov5640_reg[(209*24)+1*8+:8], w_ov5640_reg[(209*24)+2*8+:8]}	= 24'h303511;
assign	{w_ov5640_reg[(210*24)+0*8+:8], w_ov5640_reg[(210*24)+1*8+:8], w_ov5640_reg[(210*24)+2*8+:8]}	= 24'h30365D;
assign	{w_ov5640_reg[(211*24)+0*8+:8], w_ov5640_reg[(211*24)+1*8+:8], w_ov5640_reg[(211*24)+2*8+:8]}	= 24'h3c0707;
assign	{w_ov5640_reg[(212*24)+0*8+:8], w_ov5640_reg[(212*24)+1*8+:8], w_ov5640_reg[(212*24)+2*8+:8]}	= 24'h382047;
assign	{w_ov5640_reg[(213*24)+0*8+:8], w_ov5640_reg[(213*24)+1*8+:8], w_ov5640_reg[(213*24)+2*8+:8]}	= 24'h382107;
assign	{w_ov5640_reg[(214*24)+0*8+:8], w_ov5640_reg[(214*24)+1*8+:8], w_ov5640_reg[(214*24)+2*8+:8]}	= 24'h381431;
assign	{w_ov5640_reg[(215*24)+0*8+:8], w_ov5640_reg[(215*24)+1*8+:8], w_ov5640_reg[(215*24)+2*8+:8]}	= 24'h381531;
assign	{w_ov5640_reg[(216*24)+0*8+:8], w_ov5640_reg[(216*24)+1*8+:8], w_ov5640_reg[(216*24)+2*8+:8]}	= 24'h380000;
assign	{w_ov5640_reg[(217*24)+0*8+:8], w_ov5640_reg[(217*24)+1*8+:8], w_ov5640_reg[(217*24)+2*8+:8]}	= 24'h380100;
assign	{w_ov5640_reg[(218*24)+0*8+:8], w_ov5640_reg[(218*24)+1*8+:8], w_ov5640_reg[(218*24)+2*8+:8]}	= 24'h380200;
assign	{w_ov5640_reg[(219*24)+0*8+:8], w_ov5640_reg[(219*24)+1*8+:8], w_ov5640_reg[(219*24)+2*8+:8]}	= 24'h3803fa;
assign	{w_ov5640_reg[(220*24)+0*8+:8], w_ov5640_reg[(220*24)+1*8+:8], w_ov5640_reg[(220*24)+2*8+:8]}	= 24'h38040a;
assign	{w_ov5640_reg[(221*24)+0*8+:8], w_ov5640_reg[(221*24)+1*8+:8], w_ov5640_reg[(221*24)+2*8+:8]}	= 24'h38053f;
assign	{w_ov5640_reg[(222*24)+0*8+:8], w_ov5640_reg[(222*24)+1*8+:8], w_ov5640_reg[(222*24)+2*8+:8]}	= 24'h380606;
assign	{w_ov5640_reg[(223*24)+0*8+:8], w_ov5640_reg[(223*24)+1*8+:8], w_ov5640_reg[(223*24)+2*8+:8]}	= 24'h3807a9;
assign	{w_ov5640_reg[(224*24)+0*8+:8], w_ov5640_reg[(224*24)+1*8+:8], w_ov5640_reg[(224*24)+2*8+:8]}	= 24'h380805;
assign	{w_ov5640_reg[(225*24)+0*8+:8], w_ov5640_reg[(225*24)+1*8+:8], w_ov5640_reg[(225*24)+2*8+:8]}	= 24'h380900;
assign	{w_ov5640_reg[(226*24)+0*8+:8], w_ov5640_reg[(226*24)+1*8+:8], w_ov5640_reg[(226*24)+2*8+:8]}	= 24'h380a02;
assign	{w_ov5640_reg[(227*24)+0*8+:8], w_ov5640_reg[(227*24)+1*8+:8], w_ov5640_reg[(227*24)+2*8+:8]}	= 24'h380bd0;
assign	{w_ov5640_reg[(228*24)+0*8+:8], w_ov5640_reg[(228*24)+1*8+:8], w_ov5640_reg[(228*24)+2*8+:8]}	= 24'h380c06;
assign	{w_ov5640_reg[(229*24)+0*8+:8], w_ov5640_reg[(229*24)+1*8+:8], w_ov5640_reg[(229*24)+2*8+:8]}	= 24'h380d72;
assign	{w_ov5640_reg[(230*24)+0*8+:8], w_ov5640_reg[(230*24)+1*8+:8], w_ov5640_reg[(230*24)+2*8+:8]}	= 24'h380e02;
assign	{w_ov5640_reg[(231*24)+0*8+:8], w_ov5640_reg[(231*24)+1*8+:8], w_ov5640_reg[(231*24)+2*8+:8]}	= 24'h380fee;
assign	{w_ov5640_reg[(232*24)+0*8+:8], w_ov5640_reg[(232*24)+1*8+:8], w_ov5640_reg[(232*24)+2*8+:8]}	= 24'h381302;
assign	{w_ov5640_reg[(233*24)+0*8+:8], w_ov5640_reg[(233*24)+1*8+:8], w_ov5640_reg[(233*24)+2*8+:8]}	= 24'h361800;
assign	{w_ov5640_reg[(234*24)+0*8+:8], w_ov5640_reg[(234*24)+1*8+:8], w_ov5640_reg[(234*24)+2*8+:8]}	= 24'h361229;
assign	{w_ov5640_reg[(235*24)+0*8+:8], w_ov5640_reg[(235*24)+1*8+:8], w_ov5640_reg[(235*24)+2*8+:8]}	= 24'h370952;
assign	{w_ov5640_reg[(236*24)+0*8+:8], w_ov5640_reg[(236*24)+1*8+:8], w_ov5640_reg[(236*24)+2*8+:8]}	= 24'h370c03;
assign	{w_ov5640_reg[(237*24)+0*8+:8], w_ov5640_reg[(237*24)+1*8+:8], w_ov5640_reg[(237*24)+2*8+:8]}	= 24'h3a0202;
assign	{w_ov5640_reg[(238*24)+0*8+:8], w_ov5640_reg[(238*24)+1*8+:8], w_ov5640_reg[(238*24)+2*8+:8]}	= 24'h3a03e0;
assign	{w_ov5640_reg[(239*24)+0*8+:8], w_ov5640_reg[(239*24)+1*8+:8], w_ov5640_reg[(239*24)+2*8+:8]}	= 24'h3a0800;
assign	{w_ov5640_reg[(240*24)+0*8+:8], w_ov5640_reg[(240*24)+1*8+:8], w_ov5640_reg[(240*24)+2*8+:8]}	= 24'h3a096f;
assign	{w_ov5640_reg[(241*24)+0*8+:8], w_ov5640_reg[(241*24)+1*8+:8], w_ov5640_reg[(241*24)+2*8+:8]}	= 24'h3a0a00;
assign	{w_ov5640_reg[(242*24)+0*8+:8], w_ov5640_reg[(242*24)+1*8+:8], w_ov5640_reg[(242*24)+2*8+:8]}	= 24'h3a0b5c;
assign	{w_ov5640_reg[(243*24)+0*8+:8], w_ov5640_reg[(243*24)+1*8+:8], w_ov5640_reg[(243*24)+2*8+:8]}	= 24'h3a0e06;
assign	{w_ov5640_reg[(244*24)+0*8+:8], w_ov5640_reg[(244*24)+1*8+:8], w_ov5640_reg[(244*24)+2*8+:8]}	= 24'h3a0d08;
assign	{w_ov5640_reg[(245*24)+0*8+:8], w_ov5640_reg[(245*24)+1*8+:8], w_ov5640_reg[(245*24)+2*8+:8]}	= 24'h3a1402;
assign	{w_ov5640_reg[(246*24)+0*8+:8], w_ov5640_reg[(246*24)+1*8+:8], w_ov5640_reg[(246*24)+2*8+:8]}	= 24'h3a15e0;
assign	{w_ov5640_reg[(247*24)+0*8+:8], w_ov5640_reg[(247*24)+1*8+:8], w_ov5640_reg[(247*24)+2*8+:8]}	= 24'h400402;
assign	{w_ov5640_reg[(248*24)+0*8+:8], w_ov5640_reg[(248*24)+1*8+:8], w_ov5640_reg[(248*24)+2*8+:8]}	= 24'h30021c;
assign	{w_ov5640_reg[(249*24)+0*8+:8], w_ov5640_reg[(249*24)+1*8+:8], w_ov5640_reg[(249*24)+2*8+:8]}	= 24'h3006c3;
assign	{w_ov5640_reg[(250*24)+0*8+:8], w_ov5640_reg[(250*24)+1*8+:8], w_ov5640_reg[(250*24)+2*8+:8]}	= 24'h471303;
assign	{w_ov5640_reg[(251*24)+0*8+:8], w_ov5640_reg[(251*24)+1*8+:8], w_ov5640_reg[(251*24)+2*8+:8]}	= 24'h440704;
assign	{w_ov5640_reg[(252*24)+0*8+:8], w_ov5640_reg[(252*24)+1*8+:8], w_ov5640_reg[(252*24)+2*8+:8]}	= 24'h460b37;
assign	{w_ov5640_reg[(253*24)+0*8+:8], w_ov5640_reg[(253*24)+1*8+:8], w_ov5640_reg[(253*24)+2*8+:8]}	= 24'h460c20;
assign	{w_ov5640_reg[(254*24)+0*8+:8], w_ov5640_reg[(254*24)+1*8+:8], w_ov5640_reg[(254*24)+2*8+:8]}	= 24'h483716;
assign	{w_ov5640_reg[(255*24)+0*8+:8], w_ov5640_reg[(255*24)+1*8+:8], w_ov5640_reg[(255*24)+2*8+:8]}	= 24'h382404;
assign	{w_ov5640_reg[(256*24)+0*8+:8], w_ov5640_reg[(256*24)+1*8+:8], w_ov5640_reg[(256*24)+2*8+:8]}	= 24'h500183;
assign	{w_ov5640_reg[(257*24)+0*8+:8], w_ov5640_reg[(257*24)+1*8+:8], w_ov5640_reg[(257*24)+2*8+:8]}	= 24'h350300;
assign	{w_ov5640_reg[(258*24)+0*8+:8], w_ov5640_reg[(258*24)+1*8+:8], w_ov5640_reg[(258*24)+2*8+:8]}	= 24'h301602;
assign	{w_ov5640_reg[(259*24)+0*8+:8], w_ov5640_reg[(259*24)+1*8+:8], w_ov5640_reg[(259*24)+2*8+:8]}	= 24'h3b070a;
assign	{w_ov5640_reg[(260*24)+0*8+:8], w_ov5640_reg[(260*24)+1*8+:8], w_ov5640_reg[(260*24)+2*8+:8]}	= 24'h503d00;
assign	{w_ov5640_reg[(261*24)+0*8+:8], w_ov5640_reg[(261*24)+1*8+:8], w_ov5640_reg[(261*24)+2*8+:8]}	= 24'h474100;
assign	{w_ov5640_reg[(262*24)+0*8+:8], w_ov5640_reg[(262*24)+1*8+:8], w_ov5640_reg[(262*24)+2*8+:8]}	= 24'h470905;
assign	w_ov5640_reg[8191:263*24]	= {848{1'b0}};

assign	o_data	= w_ov5640_reg[i_addr*8+:8];

endmodule
